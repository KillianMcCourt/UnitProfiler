--------------------------------------------------------------------------------
--                 FixRealKCM_Freq300_uid58_T0_Freq300_uid61
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid58_T0_Freq300_uid61 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(80 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid58_T0_Freq300_uid61 is
signal Y0 :  std_logic_vector(80 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(80 downto 0);
begin
   with X  select  Y0 <= 
      "000000000000000000000000000000000000000000000000000000000000000000000000000000000" when "00000",
      "000001011000101110010000101111111011111010001110011110111100110101011110010011110" when "00001",
      "000010110001011100100001011111110111110100011100111101111001101010111100100111100" when "00010",
      "000100001010001010110010001111110011101110101011011100110110100000011010111011011" when "00011",
      "000101100010111001000010111111101111101000111001111011110011010101111001001111001" when "00100",
      "000110111011100111010011101111101011100011001000011010110000001011010111100010111" when "00101",
      "001000010100010101100100011111100111011101010110111001101101000000110101110110101" when "00110",
      "001001101101000011110101001111100011010111100101011000101001110110010100001010100" when "00111",
      "001011000101110010000101111111011111010001110011110111100110101011110010011110010" when "01000",
      "001100011110100000010110101111011011001100000010010110100011100001010000110010000" when "01001",
      "001101110111001110100111011111010111000110010000110101100000010110101111000101110" when "01010",
      "001111001111111100111000001111010011000000011111010100011101001100001101011001101" when "01011",
      "010000101000101011001000111111001110111010101101110011011010000001101011101101011" when "01100",
      "010010000001011001011001101111001010110100111100010010010110110111001010000001001" when "01101",
      "010011011010000111101010011111000110101111001010110001010011101100101000010100111" when "01110",
      "010100110010110101111011001111000010101001011001010000010000100010000110101000101" when "01111",
      "010110001011100100001011111110111110100011100111101111001101010111100100111100100" when "10000",
      "010111100100010010011100101110111010011101110110001110001010001101000011010000010" when "10001",
      "011000111101000000101101011110110110011000000100101101000111000010100001100100000" when "10010",
      "011010010101101110111110001110110010010010010011001100000011110111111111110111110" when "10011",
      "011011101110011101001110111110101110001100100001101011000000101101011110001011101" when "10100",
      "011101000111001011011111101110101010000110110000001001111101100010111100011111011" when "10101",
      "011110011111111001110000011110100110000000111110101000111010011000011010110011001" when "10110",
      "011111111000101000000001001110100001111011001101000111110111001101111001000110111" when "10111",
      "100001010001010110010001111110011101110101011011100110110100000011010111011010110" when "11000",
      "100010101010000100100010101110011001101111101010000101110000111000110101101110100" when "11001",
      "100100000010110010110011011110010101101001111000100100101101101110010100000010010" when "11010",
      "100101011011100001000100001110010001100100000111000011101010100011110010010110000" when "11011",
      "100110110100001111010100111110001101011110010101100010100111011001010000101001110" when "11100",
      "101000001100111101100101101110001001011000100100000001100100001110101110111101101" when "11101",
      "101001100101101011110110011110000101010010110010100000100001000100001101010001011" when "11110",
      "101010111110011010000111001110000001001101000000111111011101111001101011100101001" when "11111",
      "---------------------------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq300_uid58_T1_Freq300_uid64
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid58_T1_Freq300_uid64 is
    port (X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(75 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid58_T1_Freq300_uid64 is
signal Y0 :  std_logic_vector(75 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(75 downto 0);
begin
   with X  select  Y0 <= 
      "0000000000000000000000000000000000000000000000000000000000000000000000000000" when "000000",
      "0000001011000101110010000101111111011111010001110011110111100110101011110010" when "000001",
      "0000010110001011100100001011111110111110100011100111101111001101010111100101" when "000010",
      "0000100001010001010110010001111110011101110101011011100110110100000011010111" when "000011",
      "0000101100010111001000010111111101111101000111001111011110011010101111001010" when "000100",
      "0000110111011100111010011101111101011100011001000011010110000001011010111100" when "000101",
      "0001000010100010101100100011111100111011101010110111001101101000000110101111" when "000110",
      "0001001101101000011110101001111100011010111100101011000101001110110010100001" when "000111",
      "0001011000101110010000101111111011111010001110011110111100110101011110010100" when "001000",
      "0001100011110100000010110101111011011001100000010010110100011100001010000110" when "001001",
      "0001101110111001110100111011111010111000110010000110101100000010110101111001" when "001010",
      "0001111001111111100111000001111010011000000011111010100011101001100001101011" when "001011",
      "0010000101000101011001000111111001110111010101101110011011010000001101011110" when "001100",
      "0010010000001011001011001101111001010110100111100010010010110110111001010000" when "001101",
      "0010011011010000111101010011111000110101111001010110001010011101100101000011" when "001110",
      "0010100110010110101111011001111000010101001011001010000010000100010000110101" when "001111",
      "0010110001011100100001011111110111110100011100111101111001101010111100101000" when "010000",
      "0010111100100010010011100101110111010011101110110001110001010001101000011010" when "010001",
      "0011000111101000000101101011110110110011000000100101101000111000010100001101" when "010010",
      "0011010010101101110111110001110110010010010010011001100000011110111111111111" when "010011",
      "0011011101110011101001110111110101110001100100001101011000000101101011110001" when "010100",
      "0011101000111001011011111101110101010000110110000001001111101100010111100100" when "010101",
      "0011110011111111001110000011110100110000000111110101000111010011000011010110" when "010110",
      "0011111111000101000000001001110100001111011001101000111110111001101111001001" when "010111",
      "0100001010001010110010001111110011101110101011011100110110100000011010111011" when "011000",
      "0100010101010000100100010101110011001101111101010000101110000111000110101110" when "011001",
      "0100100000010110010110011011110010101101001111000100100101101101110010100000" when "011010",
      "0100101011011100001000100001110010001100100000111000011101010100011110010011" when "011011",
      "0100110110100001111010100111110001101011110010101100010100111011001010000101" when "011100",
      "0101000001100111101100101101110001001011000100100000001100100001110101111000" when "011101",
      "0101001100101101011110110011110000101010010110010100000100001000100001101010" when "011110",
      "0101010111110011010000111001110000001001101000000111111011101111001101011101" when "011111",
      "0101100010111001000010111111101111101000111001111011110011010101111001001111" when "100000",
      "0101101101111110110101000101101111001000001011101111101010111100100101000010" when "100001",
      "0101111001000100100111001011101110100111011101100011100010100011010000110100" when "100010",
      "0110000100001010011001010001101110000110101111010111011010001001111100100111" when "100011",
      "0110001111010000001011010111101101100110000001001011010001110000101000011001" when "100100",
      "0110011010010101111101011101101101000101010010111111001001010111010100001011" when "100101",
      "0110100101011011101111100011101100100100100100110011000000111101111111111110" when "100110",
      "0110110000100001100001101001101100000011110110100110111000100100101011110000" when "100111",
      "0110111011100111010011101111101011100011001000011010110000001011010111100011" when "101000",
      "0111000110101101000101110101101011000010011010001110100111110010000011010101" when "101001",
      "0111010001110010110111111011101010100001101100000010011111011000101111001000" when "101010",
      "0111011100111000101010000001101010000000111101110110010110111111011010111010" when "101011",
      "0111100111111110011100000111101001100000001111101010001110100110000110101101" when "101100",
      "0111110011000100001110001101101000111111100001011110000110001100110010011111" when "101101",
      "0111111110001010000000010011101000011110110011010001111101110011011110010010" when "101110",
      "1000001001001111110010011001100111111110000101000101110101011010001010000100" when "101111",
      "1000010100010101100100011111100111011101010110111001101101000000110101110111" when "110000",
      "1000011111011011010110100101100110111100101000101101100100100111100001101001" when "110001",
      "1000101010100001001000101011100110011011111010100001011100001110001101011100" when "110010",
      "1000110101100110111010110001100101111011001100010101010011110100111001001110" when "110011",
      "1001000000101100101100110111100101011010011110001001001011011011100101000001" when "110100",
      "1001001011110010011110111101100100111001101111111101000011000010010000110011" when "110101",
      "1001010110111000010001000011100100011001000001110000111010101000111100100110" when "110110",
      "1001100001111110000011001001100011111000010011100100110010001111101000011000" when "110111",
      "1001101101000011110101001111100011010111100101011000101001110110010100001010" when "111000",
      "1001111000001001100111010101100010110110110111001100100001011100111111111101" when "111001",
      "1010000011001111011001011011100010010110001001000000011001000011101011101111" when "111010",
      "1010001110010101001011100001100001110101011010110100010000101010010111100010" when "111011",
      "1010011001011010111101100111100001010100101100101000001000010001000011010100" when "111100",
      "1010100100100000101111101101100000110011111110011011111111110111101111000111" when "111101",
      "1010101111100110100001110011100000010011010000001111110111011110011010111001" when "111110",
      "1010111010101100010011111001011111110010100010000011101111000101000110101100" when "111111",
      "----------------------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid100
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid100 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid100 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid107
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid107 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid107 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid112
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid112 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid112 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid121
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid121 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid121 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid126
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid126 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid126 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid133
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid133 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid133 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid138
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid143
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid143 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid143 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid150
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid150 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid150 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid155
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid155 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid155 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid160
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid160 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid160 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid165
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid165 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid165 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid180
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid180 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid180 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid189
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid189 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid189 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid196
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid196 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid196 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid201
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid201 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid201 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid208
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid208 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid208 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid213
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid213 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid213 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid218
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid227
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid227 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid227 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid232
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid232 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid232 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid237
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid237 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid237 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid244
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid244 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid244 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid249
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid249 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid249 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid254
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid254 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid254 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid259
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid259 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid259 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid266
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid266 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid266 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid271
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid271 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid271 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid276
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid276 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid276 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid281
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid281 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid281 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid286
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid286 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid286 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid293
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid293 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid293 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid298
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid298 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid298 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid303
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid303 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid303 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid308
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid308 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid308 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid313
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid313 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid313 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid320
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid320 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid320 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid325
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid325 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid325 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid330
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid330 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid330 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid335
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid335 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid335 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid340
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid340 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid340 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid355
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid355 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid355 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid360
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid360 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid360 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid365
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid365 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid365 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid370
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid370 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid370 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid375
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid375 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid375 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid380
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid380 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid380 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid385
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid385 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid385 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid390
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid390 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid390 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid395
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid395 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid395 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid400
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid400 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid400 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid405
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid405 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid405 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid410
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid410 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid410 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid425
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid425 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid425 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid430
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid430 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid430 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid435
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid435 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid435 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid440
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid440 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid440 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid445
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid445 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid445 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid450
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid450 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid450 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid455
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid455 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid455 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid460
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid460 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid460 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid465
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid465 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid465 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid470
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid470 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid470 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid475
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid475 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid475 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid480
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid480 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid480 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid495
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid495 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid495 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid500
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid500 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid500 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid505
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid505 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid505 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid510
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid510 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid510 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid515
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid515 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid515 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid520
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid520 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid520 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid525
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid525 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid525 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid530
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid530 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid530 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid535
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid535 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid535 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid540
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid540 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid540 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid545
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid545 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid545 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid550
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid550 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid550 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid565
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid565 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid565 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid570
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid570 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid570 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid575
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid575 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid575 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid580
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid580 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid580 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid585
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid585 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid585 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid592
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid592 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid592 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid597
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid597 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid597 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid602
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid602 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid602 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid607
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid607 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid607 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid612
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid612 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid612 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid616
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid616 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid616 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq300_uid626
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid626 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid626 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid650
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid650 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid650 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid712
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid712 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid712 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid958
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid958 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid958 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--               FixRealKCM_Freq300_uid1483_T0_Freq300_uid1486
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1483_T0_Freq300_uid1486 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1483_T0_Freq300_uid1486 is
signal Y0 :  std_logic_vector(14 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(14 downto 0);
begin
   with X  select  Y0 <= 
      "000000000001000" when "00000",
      "000001011101011" when "00001",
      "000010111001101" when "00010",
      "000100010110000" when "00011",
      "000101110010011" when "00100",
      "000111001110101" when "00101",
      "001000101011000" when "00110",
      "001010000111011" when "00111",
      "001011100011101" when "01000",
      "001101000000000" when "01001",
      "001110011100011" when "01010",
      "001111111000101" when "01011",
      "010001010101000" when "01100",
      "010010110001011" when "01101",
      "010100001101101" when "01110",
      "010101101010000" when "01111",
      "010111000110011" when "10000",
      "011000100010101" when "10001",
      "011001111111000" when "10010",
      "011011011011011" when "10011",
      "011100110111101" when "10100",
      "011110010100000" when "10101",
      "011111110000011" when "10110",
      "100001001100101" when "10111",
      "100010101001000" when "11000",
      "100100000101010" when "11001",
      "100101100001101" when "11010",
      "100110111110000" when "11011",
      "101000011010010" when "11100",
      "101001110110101" when "11101",
      "101011010011000" when "11110",
      "101100101111010" when "11111",
      "---------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--               FixRealKCM_Freq300_uid1483_T1_Freq300_uid1489
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1483_T1_Freq300_uid1489 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1483_T1_Freq300_uid1489 is
signal Y0 :  std_logic_vector(9 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(9 downto 0);
begin
   with X  select  Y0 <= 
      "0000000000" when "00000",
      "0000010111" when "00001",
      "0000101110" when "00010",
      "0001000101" when "00011",
      "0001011100" when "00100",
      "0001110011" when "00101",
      "0010001010" when "00110",
      "0010100010" when "00111",
      "0010111001" when "01000",
      "0011010000" when "01001",
      "0011100111" when "01010",
      "0011111110" when "01011",
      "0100010101" when "01100",
      "0100101100" when "01101",
      "0101000011" when "01110",
      "0101011010" when "01111",
      "0101110001" when "10000",
      "0110001000" when "10001",
      "0110011111" when "10010",
      "0110110111" when "10011",
      "0111001110" when "10100",
      "0111100101" when "10101",
      "0111111100" when "10110",
      "1000010011" when "10111",
      "1000101010" when "11000",
      "1001000001" when "11001",
      "1001011000" when "11010",
      "1001101111" when "11011",
      "1010000110" when "11100",
      "1010011101" when "11101",
      "1010110100" when "11110",
      "1011001100" when "11111",
      "----------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--               FixRealKCM_Freq300_uid1483_T2_Freq300_uid1492
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1483_T2_Freq300_uid1492 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1483_T2_Freq300_uid1492 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "000",
      "00011" when "001",
      "00110" when "010",
      "01001" when "011",
      "01100" when "100",
      "01110" when "101",
      "10001" when "110",
      "10100" when "111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_23_3_Freq300_uid1496
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid1496 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid1496 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--               FixRealKCM_Freq300_uid1510_T0_Freq300_uid1513
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1510_T0_Freq300_uid1513 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(66 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1510_T0_Freq300_uid1513 is
signal Y0 :  std_logic_vector(66 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(66 downto 0);
begin
   with X  select  Y0 <= 
      "0000000000000000000000000000000000000000000000000000000000000000000" when "00000",
      "0000010110001011100100001011111110111110100011100111101111001101011" when "00001",
      "0000101100010111001000010111111101111101000111001111011110011010110" when "00010",
      "0001000010100010101100100011111100111011101010110111001101101000001" when "00011",
      "0001011000101110010000101111111011111010001110011110111100110101100" when "00100",
      "0001101110111001110100111011111010111000110010000110101100000010111" when "00101",
      "0010000101000101011001000111111001110111010101101110011011010000010" when "00110",
      "0010011011010000111101010011111000110101111001010110001010011101101" when "00111",
      "0010110001011100100001011111110111110100011100111101111001101011000" when "01000",
      "0011000111101000000101101011110110110011000000100101101000111000011" when "01001",
      "0011011101110011101001110111110101110001100100001101011000000101101" when "01010",
      "0011110011111111001110000011110100110000000111110101000111010011000" when "01011",
      "0100001010001010110010001111110011101110101011011100110110100000011" when "01100",
      "0100100000010110010110011011110010101101001111000100100101101101110" when "01101",
      "0100110110100001111010100111110001101011110010101100010100111011001" when "01110",
      "0101001100101101011110110011110000101010010110010100000100001000100" when "01111",
      "0101100010111001000010111111101111101000111001111011110011010101111" when "10000",
      "0101111001000100100111001011101110100111011101100011100010100011010" when "10001",
      "0110001111010000001011010111101101100110000001001011010001110000101" when "10010",
      "0110100101011011101111100011101100100100100100110011000000111110000" when "10011",
      "0110111011100111010011101111101011100011001000011010110000001011011" when "10100",
      "0111010001110010110111111011101010100001101100000010011111011000110" when "10101",
      "0111100111111110011100000111101001100000001111101010001110100110001" when "10110",
      "0111111110001010000000010011101000011110110011010001111101110011100" when "10111",
      "1000010100010101100100011111100111011101010110111001101101000000111" when "11000",
      "1000101010100001001000101011100110011011111010100001011100001110010" when "11001",
      "1001000000101100101100110111100101011010011110001001001011011011101" when "11010",
      "1001010110111000010001000011100100011001000001110000111010101001000" when "11011",
      "1001101101000011110101001111100011010111100101011000101001110110011" when "11100",
      "1010000011001111011001011011100010010110001001000000011001000011101" when "11101",
      "1010011001011010111101100111100001010100101100101000001000010001000" when "11110",
      "1010101111100110100001110011100000010011010000001111110111011110011" when "11111",
      "-------------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--               FixRealKCM_Freq300_uid1510_T1_Freq300_uid1516
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1510_T1_Freq300_uid1516 is
    port (X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1510_T1_Freq300_uid1516 is
signal Y0 :  std_logic_vector(61 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(61 downto 0);
begin
   with X  select  Y0 <= 
      "00000000000000000000000000000000000000000000000000000000000000" when "000000",
      "00000010110001011100100001011111110111110100011100111101111010" when "000001",
      "00000101100010111001000010111111101111101000111001111011110011" when "000010",
      "00001000010100010101100100011111100111011101010110111001101101" when "000011",
      "00001011000101110010000101111111011111010001110011110111100111" when "000100",
      "00001101110111001110100111011111010111000110010000110101100000" when "000101",
      "00010000101000101011001000111111001110111010101101110011011010" when "000110",
      "00010011011010000111101010011111000110101111001010110001010100" when "000111",
      "00010110001011100100001011111110111110100011100111101111001101" when "001000",
      "00011000111101000000101101011110110110011000000100101101000111" when "001001",
      "00011011101110011101001110111110101110001100100001101011000001" when "001010",
      "00011110011111111001110000011110100110000000111110101000111010" when "001011",
      "00100001010001010110010001111110011101110101011011100110110100" when "001100",
      "00100100000010110010110011011110010101101001111000100100101110" when "001101",
      "00100110110100001111010100111110001101011110010101100010100111" when "001110",
      "00101001100101101011110110011110000101010010110010100000100001" when "001111",
      "00101100010111001000010111111101111101000111001111011110011011" when "010000",
      "00101111001000100100111001011101110100111011101100011100010100" when "010001",
      "00110001111010000001011010111101101100110000001001011010001110" when "010010",
      "00110100101011011101111100011101100100100100100110011000001000" when "010011",
      "00110111011100111010011101111101011100011001000011010110000001" when "010100",
      "00111010001110010110111111011101010100001101100000010011111011" when "010101",
      "00111100111111110011100000111101001100000001111101010001110101" when "010110",
      "00111111110001010000000010011101000011110110011010001111101110" when "010111",
      "01000010100010101100100011111100111011101010110111001101101000" when "011000",
      "01000101010100001001000101011100110011011111010100001011100010" when "011001",
      "01001000000101100101100110111100101011010011110001001001011011" when "011010",
      "01001010110111000010001000011100100011001000001110000111010101" when "011011",
      "01001101101000011110101001111100011010111100101011000101001111" when "011100",
      "01010000011001111011001011011100010010110001001000000011001000" when "011101",
      "01010011001011010111101100111100001010100101100101000001000010" when "011110",
      "01010101111100110100001110011100000010011010000001111110111100" when "011111",
      "01011000101110010000101111111011111010001110011110111100110101" when "100000",
      "01011011011111101101010001011011110010000010111011111010101111" when "100001",
      "01011110010001001001110010111011101001110111011000111000101001" when "100010",
      "01100001000010100110010100011011100001101011110101110110100010" when "100011",
      "01100011110100000010110101111011011001100000010010110100011100" when "100100",
      "01100110100101011111010111011011010001010100101111110010010110" when "100101",
      "01101001010110111011111000111011001001001001001100110000001111" when "100110",
      "01101100001000011000011010011011000000111101101001101110001001" when "100111",
      "01101110111001110100111011111010111000110010000110101100000011" when "101000",
      "01110001101011010001011101011010110000100110100011101001111101" when "101001",
      "01110100011100101101111110111010101000011011000000100111110110" when "101010",
      "01110111001110001010100000011010100000001111011101100101110000" when "101011",
      "01111001111111100111000001111010011000000011111010100011101010" when "101100",
      "01111100110001000011100011011010001111111000010111100001100011" when "101101",
      "01111111100010100000000100111010000111101100110100011111011101" when "101110",
      "10000010010011111100100110011001111111100001010001011101010111" when "101111",
      "10000101000101011001000111111001110111010101101110011011010000" when "110000",
      "10000111110110110101101001011001101111001010001011011001001010" when "110001",
      "10001010101000010010001010111001100110111110101000010111000100" when "110010",
      "10001101011001101110101100011001011110110011000101010100111101" when "110011",
      "10010000001011001011001101111001010110100111100010010010110111" when "110100",
      "10010010111100100111101111011001001110011011111111010000110001" when "110101",
      "10010101101110000100010000111001000110010000011100001110101010" when "110110",
      "10011000011111100000110010011000111110000100111001001100100100" when "110111",
      "10011011010000111101010011111000110101111001010110001010011110" when "111000",
      "10011110000010011001110101011000101101101101110011001000010111" when "111001",
      "10100000110011110110010110111000100101100010010000000110010001" when "111010",
      "10100011100101010010111000011000011101010110101101000100001011" when "111011",
      "10100110010110101111011001111000010101001011001010000010000100" when "111100",
      "10101001001000001011111011011000001100111111100110111111111110" when "111101",
      "10101011111001101000011100111000000100110100000011111101111000" when "111110",
      "10101110101011000100111110010111111100101000100000111011110001" when "111111",
      "--------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--        compressedTable_Freq300_uid1527_subsampling_Freq300_uid1529
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq300_uid1527_subsampling_Freq300_uid1529 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of compressedTable_Freq300_uid1527_subsampling_Freq300_uid1529 is
signal Y0 :  std_logic_vector(8 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(8 downto 0);
begin
   with X  select  Y0 <= 
      "100000000" when "0000000",
      "100000010" when "0000001",
      "100000100" when "0000010",
      "100000110" when "0000011",
      "100001000" when "0000100",
      "100001010" when "0000101",
      "100001100" when "0000110",
      "100001110" when "0000111",
      "100010000" when "0001000",
      "100010010" when "0001001",
      "100010100" when "0001010",
      "100010110" when "0001011",
      "100011001" when "0001100",
      "100011011" when "0001101",
      "100011101" when "0001110",
      "100011111" when "0001111",
      "100100010" when "0010000",
      "100100100" when "0010001",
      "100100110" when "0010010",
      "100101000" when "0010011",
      "100101011" when "0010100",
      "100101101" when "0010101",
      "100110000" when "0010110",
      "100110010" when "0010111",
      "100110100" when "0011000",
      "100110111" when "0011001",
      "100111001" when "0011010",
      "100111100" when "0011011",
      "100111110" when "0011100",
      "101000001" when "0011101",
      "101000011" when "0011110",
      "101000110" when "0011111",
      "101001000" when "0100000",
      "101001011" when "0100001",
      "101001101" when "0100010",
      "101010000" when "0100011",
      "101010011" when "0100100",
      "101010101" when "0100101",
      "101011000" when "0100110",
      "101011011" when "0100111",
      "101011101" when "0101000",
      "101100000" when "0101001",
      "101100011" when "0101010",
      "101100110" when "0101011",
      "101101001" when "0101100",
      "101101011" when "0101101",
      "101101110" when "0101110",
      "101110001" when "0101111",
      "101110100" when "0110000",
      "101110111" when "0110001",
      "101111010" when "0110010",
      "101111101" when "0110011",
      "110000000" when "0110100",
      "110000011" when "0110101",
      "110000110" when "0110110",
      "110001001" when "0110111",
      "110001100" when "0111000",
      "110001111" when "0111001",
      "110010010" when "0111010",
      "110010101" when "0111011",
      "110011001" when "0111100",
      "110011100" when "0111101",
      "110011111" when "0111110",
      "110100010" when "0111111",
      "010011011" when "1000000",
      "010011100" when "1000001",
      "010011101" when "1000010",
      "010011110" when "1000011",
      "010100000" when "1000100",
      "010100001" when "1000101",
      "010100010" when "1000110",
      "010100011" when "1000111",
      "010100101" when "1001000",
      "010100110" when "1001001",
      "010100111" when "1001010",
      "010101001" when "1001011",
      "010101010" when "1001100",
      "010101011" when "1001101",
      "010101101" when "1001110",
      "010101110" when "1001111",
      "010101111" when "1010000",
      "010110001" when "1010001",
      "010110010" when "1010010",
      "010110100" when "1010011",
      "010110101" when "1010100",
      "010110110" when "1010101",
      "010111000" when "1010110",
      "010111001" when "1010111",
      "010111011" when "1011000",
      "010111100" when "1011001",
      "010111110" when "1011010",
      "010111111" when "1011011",
      "011000001" when "1011100",
      "011000010" when "1011101",
      "011000100" when "1011110",
      "011000101" when "1011111",
      "011000111" when "1100000",
      "011001000" when "1100001",
      "011001010" when "1100010",
      "011001100" when "1100011",
      "011001101" when "1100100",
      "011001111" when "1100101",
      "011010000" when "1100110",
      "011010010" when "1100111",
      "011010100" when "1101000",
      "011010101" when "1101001",
      "011010111" when "1101010",
      "011011001" when "1101011",
      "011011010" when "1101100",
      "011011100" when "1101101",
      "011011110" when "1101110",
      "011100000" when "1101111",
      "011100001" when "1110000",
      "011100011" when "1110001",
      "011100101" when "1110010",
      "011100111" when "1110011",
      "011101001" when "1110100",
      "011101010" when "1110101",
      "011101100" when "1110110",
      "011101110" when "1110111",
      "011110000" when "1111000",
      "011110010" when "1111001",
      "011110100" when "1111010",
      "011110110" when "1111011",
      "011111000" when "1111100",
      "011111010" when "1111101",
      "011111100" when "1111110",
      "011111110" when "1111111",
      "---------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         coeffTable_Freq300_uid1536
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity coeffTable_Freq300_uid1536 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(94 downto 0)   );
end entity;

architecture arch of coeffTable_Freq300_uid1536 is
signal Y0 :  std_logic_vector(94 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(94 downto 0);
begin
   with X  select  Y0 <= 
      "00000000000000010000000000000000001001100000001000000000000000000101000100000000000000000100000" when "0000000",
      "00000000000010010000000000000010010100000000011000000000000000100101000100000000000000001100000" when "0000001",
      "00000000000110010000000000001010011110100000101000000000000001100101000100000000000000010100000" when "0000010",
      "00000000001100010000000000011100101001100000111000000000000011000101000100000000000000011100000" when "0000011",
      "00000000010100010000000000111100110100000001001000000000000101000101000100000000000000100100000" when "0000100",
      "00000000011110010000000001101110111110100001011000000000000111100101000100000000000000101100001" when "0000101",
      "00000000101010010000000010110111001001100001101000000000001010100101000100000000000000110100000" when "0000110",
      "00000000111000010000000100011001010100100001111000000000001110000101000100000000000000111011111" when "0000111",
      "00000001001000010000000110011001011111000010001000000000010010000101000100000000000001000100000" when "0001000",
      "00000001011010010000001000111011101010000010011000000000010110100101000100000000000001001100000" when "0001001",
      "00000001101110010000001100000011110101000010101000000000011011100101000100000000000001010100000" when "0001010",
      "00000010000100010000001111110110000000000010111000000000100001000101000100000000000001011100000" when "0001011",
      "00000010011100010000010100010110001011100011001000000000100111000101001100000000000001100100000" when "0001100",
      "00000010110110010000011001101000010110100011011000000000101101100101001100000000000001101100001" when "0001101",
      "00000011010010010000011111110000100010100011101000000000110100100101001100000000000001110011111" when "0001110",
      "00000011110000010000100110110010101110000011111000000000111100000101001100000000000001111100000" when "0001111",
      "00000100010000010000101110110010111010000100001000000001000100000101001100000000000010000100000" when "0010000",
      "00000100110010010000110111110101000110100100011000000001001100100101010100000000000010001100000" when "0010001",
      "00000101010110010001000001111101010011000100101000000001010101100101010100000000000010010100000" when "0010010",
      "00000101111100010001001101001111100000000100111000000001011111000101010100000000000010011011111" when "0010011",
      "00000110100100010001011001101111101101000101001000000001101001000101011100000000000010100100000" when "0010100",
      "00000111001110010001100111100001111010100101011000000001110011100101011100000000000010101100001" when "0010101",
      "00000111111010010001110110101010001001000101101000000001111110100101100100000000000010110100000" when "0010110",
      "00001000101000010010000111001100010111100101111000000010001010000101100100000000000010111100000" when "0010111",
      "00001001011000010010011001001100100110100110001000000010010110000101101100000000000011000100001" when "0011000",
      "00001010001010010010101100101110110110100110011000000010100010100101101100000000000011001100000" when "0011001",
      "00001010111110010011000001110111000111000110101000000010101111100101110100000000000011010100000" when "0011010",
      "00001011110100010011011000101001011000000110111000000010111101000101111100000000000011011100000" when "0011011",
      "00001100101100010011110001001001101001100111001000000011001011000110000100000000000011100100001" when "0011100",
      "00001101100110010100001011011011111100100111011000000011011001100110000100000000000011101100000" when "0011101",
      "00001110100010010100100111100100010000000111101000000011101000100110001100000000000011110100000" when "0011110",
      "00001111100000010101000101100110100100000111111000000011111000000110010100000000000011111100001" when "0011111",
      "00010000100000010101100101100110111001101000001000000100001000000110011100000000000100000100000" when "0100000",
      "00010001100010010110000111101001010000001000011000000100011000100110100100000000000100001100000" when "0100001",
      "00010010100110010110101011110001100111101000101000000100101001100110101100000000000100010100000" when "0100010",
      "00010011101100010111010010000100000000001000111000000100111011000110111100000000000100011100000" when "0100011",
      "00010100110100010111111010100100011010001001001000000101001101000111000100000000000100100100000" when "0100100",
      "00010101111110011000100101010110110101001001011000000101011111100111001100000000000100101100000" when "0100101",
      "00010111001010011001010010011111010001101001101000000101110010100111011100000000000100110100000" when "0100110",
      "00011000011000011010000010000001101111101001111000000110000110000111100100000000000100111100000" when "0100111",
      "00011001101000011010110100000010001111001010001000000110011010000111110100000000000101000100000" when "0101000",
      "00011010111010011011101000100100110000001010011000000110101110100111111100000000000101001100001" when "0101001",
      "00011100001110011100011111101101010011001010101000000111000011101000001100000000000101010100000" when "0101010",
      "00011101100100011101011001011111110111101010111000000111011001001000011100000000000101011100000" when "0101011",
      "00011110111100011110010110000000011110001011001000000111101111001000101100000000000101100100000" when "0101100",
      "00100000010110011111010101010011000110001011011000001000000101101000111100000000000101101100001" when "0101101",
      "00100001110010100000010111011011110000101011101000001000011100101001001100000000000101110100001" when "0101110",
      "00100011010000100001011100011110011101001011111000001000110100001001011100000000000101111100000" when "0101111",
      "00100100110000100010100100011111001011101100001000001001001100001001101100000000000110000100001" when "0110000",
      "00100110010010100011101111100001111100101100011000001001100100101001111100000000000110001100001" when "0110001",
      "00100111110110100100111101101010110000001100101000001001111101101010010100000000000110010100001" when "0110010",
      "00101001011100100110001110111101100110001100111000001010010111001010100100000000000110011100000" when "0110011",
      "00101011000100100111100011011110011110101101001000001010110001001010111100000000000110100100000" when "0110100",
      "00101100101110101000111011010001011001101101011000001011001011101011010100000000000110101100001" when "0110101",
      "00101110011010101010010110011010010111101101101000001011100110101011101100000000000110110100000" when "0110110",
      "00110000001000101011110100111101011000001101111000001100000010001100000100000000000110111100001" when "0110111",
      "00110001111000101101010110111110011100001110001000001100011110001100011100000000000111000100001" when "0111000",
      "00110011101010101110111100100001100011001110011000001100111010101100110100000000000111001100001" when "0111001",
      "00110101011110110000100101101010101101001110101000001101010111101101001100000000000111010100001" when "0111010",
      "00110111010100110010010010011101111010101110111000001101110101001101101100000000000111011100001" when "0111011",
      "00111001001100110100000010111111001011101111001000001110010011001110000100000000000111100100001" when "0111100",
      "00111011000110110101110111010010100000101111011000001110110001101110100100000000000111101100000" when "0111101",
      "00111101000010110111101111011011111000101111101000001111010000101110111100000000000111110100001" when "0111110",
      "00111111000000111001101011011111010100101111111000001111110000001111011100000000000111111100001" when "0111111",
      "01000001000000111011101011100000110100110000001000010000010000001111111100000000001000000100001" when "1000000",
      "01000011000010111101101111100100011000110000011000010000110000110000011100000000001000001100010" when "1000001",
      "01000101000110111111110111101110000001010000101000010001010001110001000100000000001000010100001" when "1000010",
      "01000111001101000010000100000001101101110000111000010001110011010001100100000000001000011100001" when "1000011",
      "01001001010101000100010100100011011110110001001000010010010101010010001100000000001000100100001" when "1000100",
      "01001011011111000110101001010111010100010001011000010010110111110010101100000000001000101100010" when "1000101",
      "01001101101011001001000010100001001110110001101000010011011010110011010100000000001000110100001" when "1000110",
      "01001111111001001011100000000101001110010001111000010011111110010011111100000000001000111100001" when "1000111",
      "01010010001001001110000010000111010010010010001000010100100010010100100100000000001001000100001" when "1001000",
      "01010100011011010000101000101011011011110010011000010101000110110101001100000000001001001100001" when "1001001",
      "01010110101111010011010011110101101010010010101000010101101011110101111100000000001001010100001" when "1001010",
      "01011001000101010110000011101001111110010010111000010110010001010110100100000000001001011100001" when "1001011",
      "01011011011101011000111000001100010111110011001000010110110111010111010100000000001001100100001" when "1001100",
      "01011101110111011011110001100000110111010011011000010111011101111000000100000000001001101100001" when "1001101",
      "01100000010011011110101111101011011100010011101000011000000100111000101100000000001001110100001" when "1001110",
      "01100010110001100001110010110000000111010011111000011000101100011001100100000000001001111100010" when "1001111",
      "01100101010001100100111010110010111000110100001000011001010100011010010100000000001010000100010" when "1010000",
      "01100111110011101000000111110111110000010100011000011001111100111011000100000000001010001100010" when "1010001",
      "01101010010111101011011010000010101110110100101000011010100101111011111100000000001010010100001" when "1010010",
      "01101100111101101110110001010111110011010100111000011011001111011100110100000000001010011100010" when "1010011",
      "01101111100101110010001101111010111111010101001000011011111001011101100100000000001010100100001" when "1010100",
      "01110010001111110101101111110000010001110101011000011100100011111110011100000000001010101100010" when "1010101",
      "01110100111011111001010110111011101011110101101000011101001110111111011100000000001010110100001" when "1010110",
      "01110111101001111101000011100001001100110101111000011101111010100000010100000000001010111100001" when "1010111",
      "01111010011010000000110101100100110101010110001000011110100110100001010100000000001011000100010" when "1011000",
      "01111101001100000100101101001010100101010110011000011111010011000010001100000000001011001100010" when "1011001",
      "10000000000000001000101010010110011101010110101000100000000000000011001100000000001011010100010" when "1011010",
      "10000010110110001100101101001100011101010110111000100000101101100100001100000000001011011100010" when "1011011",
      "10000101101110010000110101110000100101110111001000100001011011100101010100000000001011100100010" when "1011100",
      "10001000101000010101000100000110110110010111011000100010001010000110010100000000001011101100010" when "1011101",
      "10001011100100011001011000010011001111010111101000100010111001000111011100000000001011110100010" when "1011110",
      "10001110100010011101110010011001110001010111111000100011101000101000100100000000001011111100010" when "1011111",
      "10010001100010100010010010011110011011111000001000100100011000101001101100000000001100000100010" when "1100000",
      "10010100100100100110111000100101001111111000011000100101001001001010110100000000001100001100010" when "1100001",
      "10010111101000101011100100110010001100111000101000100101111010001011111100000000001100010100010" when "1100010",
      "10011010101110110000010111001001010011011000111000100110101011101101001100000000001100011100010" when "1100011",
      "10011101110110110101001111101110100011111001001000100111011101101110010100000000001100100100010" when "1100100",
      "10100001000000111010001110100101111101111001011000101000010000001111100100000000001100101100010" when "1100101",
      "10100100001100111111010011110011100001111001101000101001000011010000111100000000001100110100011" when "1100110",
      "10100111011011000100011111011011010000011001111000101001110110110010001100000000001100111100011" when "1100111",
      "10101010101011001001110001100001001001011010001000101010101010110011100100000000001101000100011" when "1101000",
      "10101101111101001111001010001001001100111010011000101011011111010100110100000000001101001100011" when "1101001",
      "10110001010001010100101001010111011011011010101000101100010100010110001100000000001101010100011" when "1101010",
      "10110100100111011010001111001111110100111010111000101101001001110111100100000000001101011100011" when "1101011",
      "10110111111111011111111011110110011001111011001000101101111111111001000100000000001101100100010" when "1101100",
      "10111011011001100101101111001111001001111011011000101110110110011010011100000000001101101100011" when "1101101",
      "10111110110101101011101001011110000101111011101000101111101101011011111100000000001101110100100" when "1101110",
      "11000010010011110001101010100111001101111011111000110000100100111101011100000000001101111100011" when "1101111",
      "11000101110011110111110010101110100010011100001000110001011100111111000100000000001110000100010" when "1110000",
      "11001001010101111110000001111000000010011100011000110010010101100000100100000000001110001100100" when "1110001",
      "11001100111010000100011000000111101111111100101000110011001110100010001100000000001110010100011" when "1110010",
      "11010000100000001010110101100001101001011100111000110100001000000011110100000000001110011100100" when "1110011",
      "11010100001000010001011010001001110000011101001000110101000010000101011100000000001110100100011" when "1110100",
      "11010111110010011000000110000100000100011101011000110101111100100111000100000000001110101100100" when "1110101",
      "11011011011110011110111001010100100110011101101000110110110111101000110100000000001110110100011" when "1110110",
      "11011111001100100101110011111111010101011101111000110111110011001010100100000000001110111100100" when "1110111",
      "11100010111100101100110110001000010010111110001000111000101111001100010100000000001111000100100" when "1111000",
      "11100110101110110011111111110011011110011110011000111001101011101110000100000000001111001100100" when "1111001",
      "11101010100010111011010001000100111000011110101000111010101000101111111100000000001111010100011" when "1111010",
      "11101110011001000010101010000000100000111110111000111011100110010001101100000000001111011100100" when "1111011",
      "11110010010001001010001010101010011000011111001000111100100100010011100100000000001111100100100" when "1111100",
      "11110110001011010001110011000110011110111111011000111101100010110101100100000000001111101100100" when "1111101",
      "11111010000111011001100011011000110100111111101000111110100001110111011100000000001111110100100" when "1111110",
      "11111110000101100001011011100101011010011111111000111111100001011001011100000000001111111100100" when "1111111",
      "-----------------------------------------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1548
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1548 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1548 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1553
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1553 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1553 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1558
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1558 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1558 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1563
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1563 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1563 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1568
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1568 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1568 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1573
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1573 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1573 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1578
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1578 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1578 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1583
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1583 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1583 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1588
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1588 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1588 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1593
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1593 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1593 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1598
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1598 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1598 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1603
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1603 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1603 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1608
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1608 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1608 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1613
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1613 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1613 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1618
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1618 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1618 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1623
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1623 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1623 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1628
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1628 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1628 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1633
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1633 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1633 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1638
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1638 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1638 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1643
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1643 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1643 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1648
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1648 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1648 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1653
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1653 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1653 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1658
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1658 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1658 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1663
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1663 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1663 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1668
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1668 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1668 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1673
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1673 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1673 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1678
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1678 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1678 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1683
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1683 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1683 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1688
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1688 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1688 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1693
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1693 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1693 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1698
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1698 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1698 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1703
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1703 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1703 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1708
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1708 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1708 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1713
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1713 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1713 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1718
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1718 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1718 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1723
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1723 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1723 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1730
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1730 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1730 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1735
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1735 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1735 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1740
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1740 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1740 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1745
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1745 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1745 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1750
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1750 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1750 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "01000" when "11000",
      "00111" when "11001",
      "00110" when "11010",
      "00101" when "11011",
      "00100" when "11100",
      "00011" when "11101",
      "00010" when "11110",
      "00001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1755
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1755 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1755 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_23_3_Freq300_uid1759
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid1759 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid1759 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid1763
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid1763 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid1763 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_14_3_Freq300_uid1767
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid1767 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid1767 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid1775
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid1775 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid1775 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid1809
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid1809 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid1809 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2022
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2022 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2022 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2027
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2027 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2027 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2032
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2032 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2032 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2037
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2037 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2037 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2042
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2042 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2042 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2047
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2047 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2047 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2052
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2052 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2052 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2057
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2057 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2057 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2062
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2062 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2062 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2067
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2067 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2067 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2072
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2072 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2072 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2077
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2077 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2077 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2082
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2082 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2082 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2087
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2087 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2087 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2092
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2092 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2092 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2097
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2097 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2097 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2102
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2102 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2102 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2107
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2107 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2107 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2112
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2112 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2112 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2117
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2117 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2117 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2122
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2122 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2122 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2127
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2127 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2127 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2132
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2132 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2132 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2137
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2137 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2137 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2142
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2142 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2142 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2147
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2147 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2147 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2152
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2152 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2152 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2157
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2157 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2157 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2162
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2162 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2162 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "01000" when "11000",
      "00111" when "11001",
      "00110" when "11010",
      "00101" when "11011",
      "00100" when "11100",
      "00011" when "11101",
      "00010" when "11110",
      "00001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2167
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2167 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2167 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2172
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2172 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2172 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2177
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2177 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2177 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2182
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2182 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2182 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2187
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2187 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2187 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2192
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2192 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2192 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2197
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2197 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2197 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2202
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2202 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2202 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2207
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2207 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2207 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2212
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2212 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2212 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2217
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2217 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2217 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2222
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2222 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2222 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2227
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2227 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2227 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2232
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2232 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2232 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2237
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2237 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2237 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2242
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2242 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2242 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2247
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2247 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2247 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2252
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2252 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2252 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_23_3_Freq300_uid2256
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid2256 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid2256 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid2264
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid2264 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid2264 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid2272
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid2272 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid2272 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_14_3_Freq300_uid2288
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid2288 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid2288 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid2314
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid2314 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid2314 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2597
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2597 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2597 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2606
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2606 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2606 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2613
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2613 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2613 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2618
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2618 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2618 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2625
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2625 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2625 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2630
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2630 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2630 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2635
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2635 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2635 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2644
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2644 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2644 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2649
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2649 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2649 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2654
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2654 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2654 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2661
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2661 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2661 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2666
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2666 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2666 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2671
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2671 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2671 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2676
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2676 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2676 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2689
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2689 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2689 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2698
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2698 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2698 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2705
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2705 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2705 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2710
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2710 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2710 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2717
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2717 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2717 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2722
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2722 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2722 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2727
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2727 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2727 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2736
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2736 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2736 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2741
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2741 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2741 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2746
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2746 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2746 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2751
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2751 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2751 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2756
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2756 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2756 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2761
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2761 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2761 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2766
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2766 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2766 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2771
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2771 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2771 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2776
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2776 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2776 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2781
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2781 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2781 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2786
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2786 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2786 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2791
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2791 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2791 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2796
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2796 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2796 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2801
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2801 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2801 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2806
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2806 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2806 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2811
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2811 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2811 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2816
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2816 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2816 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2821
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2821 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2821 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid2826
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid2826 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid2826 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_23_3_Freq300_uid2830
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid2830 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid2830 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid2834
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid2834 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid2834 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid2838
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid2838 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid2838 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_14_3_Freq300_uid2848
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid2848 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid2848 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid3032
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid3032 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid3032 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_64_Freq300_uid5
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_64_Freq300_uid5 is
    port (clk : in std_logic;
          X : in  std_logic_vector(63 downto 0);
          Y : in  std_logic_vector(63 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(63 downto 0)   );
end entity;

architecture arch of IntAdder_64_Freq300_uid5 is
signal Rtmp_c0 :  std_logic_vector(63 downto 0);
begin
   Rtmp_c0 <= X + Y + Cin;
   R <= Rtmp_c0;
end architecture;

--------------------------------------------------------------------------------
--                            LZC_52_Freq300_uid7
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: I
-- Output signals: O

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZC_52_Freq300_uid7 is
    port (clk, ce_1 : in std_logic;
          I : in  std_logic_vector(51 downto 0);
          O : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of LZC_52_Freq300_uid7 is
signal level6_c0 :  std_logic_vector(62 downto 0);
signal digit5_c0, digit5_c1 :  std_logic;
signal level5_c0 :  std_logic_vector(30 downto 0);
signal digit4_c0, digit4_c1 :  std_logic;
signal level4_c0, level4_c1 :  std_logic_vector(14 downto 0);
signal digit3_c0, digit3_c1 :  std_logic;
signal level3_c1 :  std_logic_vector(6 downto 0);
signal digit2_c1 :  std_logic;
signal level2_c1 :  std_logic_vector(2 downto 0);
signal lowBits_c1 :  std_logic_vector(1 downto 0);
signal outHighBits_c1 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               digit5_c1 <= digit5_c0;
               digit4_c1 <= digit4_c0;
               level4_c1 <= level4_c0;
               digit3_c1 <= digit3_c0;
            end if;
         end if;
      end process;
   -- pad input to the next power of two minus 1
   level6_c0 <= I & "11111111111";
   -- Main iteration for large inputs
   digit5_c0<= '1' when level6_c0(62 downto 31) = "00000000000000000000000000000000" else '0';
   level5_c0<= level6_c0(30 downto 0) when digit5_c0='1' else level6_c0(62 downto 32);
   digit4_c0<= '1' when level5_c0(30 downto 15) = "0000000000000000" else '0';
   level4_c0<= level5_c0(14 downto 0) when digit4_c0='1' else level5_c0(30 downto 16);
   digit3_c0<= '1' when level4_c0(14 downto 7) = "00000000" else '0';
   level3_c1<= level4_c1(6 downto 0) when digit3_c1='1' else level4_c1(14 downto 8);
   digit2_c1<= '1' when level3_c1(6 downto 3) = "0000" else '0';
   level2_c1<= level3_c1(2 downto 0) when digit2_c1='1' else level3_c1(6 downto 4);
   -- Finish counting with one LUT
   with level2_c1  select  lowBits_c1 <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits_c1 <= digit5_c1 & digit4_c1 & digit3_c1 & digit2_c1 & "";
   O <= outHighBits_c1 & lowBits_c1 ;
end architecture;

--------------------------------------------------------------------------------
--                           LZOC_66_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: I OZB
-- Output signals: O

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_66_Freq300_uid11 is
    port (clk, ce_1, ce_2 : in std_logic;
          I : in  std_logic_vector(65 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of LZOC_66_Freq300_uid11 is
signal sozb_c0, sozb_c1, sozb_c2 :  std_logic;
signal level7_c0 :  std_logic_vector(126 downto 0);
signal digit6_c0, digit6_c1, digit6_c2 :  std_logic;
signal level6_c0, level6_c1 :  std_logic_vector(62 downto 0);
signal digit5_c1, digit5_c2 :  std_logic;
signal level5_c1 :  std_logic_vector(30 downto 0);
signal digit4_c1, digit4_c2 :  std_logic;
signal level4_c1, level4_c2 :  std_logic_vector(14 downto 0);
signal digit3_c2 :  std_logic;
signal level3_c2 :  std_logic_vector(6 downto 0);
signal digit2_c2 :  std_logic;
signal level2_c2 :  std_logic_vector(2 downto 0);
signal z_c2 :  std_logic_vector(2 downto 0);
signal lowBits_c2 :  std_logic_vector(1 downto 0);
signal outHighBits_c2 :  std_logic_vector(4 downto 0);
signal OZB_c1, OZB_c2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sozb_c1 <= sozb_c0;
               digit6_c1 <= digit6_c0;
               level6_c1 <= level6_c0;
               OZB_c1 <= OZB;
            end if;
            if ce_2 = '1' then
               sozb_c2 <= sozb_c1;
               digit6_c2 <= digit6_c1;
               digit5_c2 <= digit5_c1;
               digit4_c2 <= digit4_c1;
               level4_c2 <= level4_c1;
               OZB_c2 <= OZB_c1;
            end if;
         end if;
      end process;
   sozb_c0 <= OZB;
   -- pad input to the next power of two minus 1
   level7_c0 <= I & (60 downto 0 => not sozb_c0);
   -- Main iteration for large inputs
   digit6_c0<= '1' when level7_c0(126 downto 63) = (63 downto 0 => sozb_c0) else '0';
   level6_c0<= level7_c0(62 downto 0) when digit6_c0='1' else level7_c0(126 downto 64);
   digit5_c1<= '1' when level6_c1(62 downto 31) = (31 downto 0 => sozb_c1) else '0';
   level5_c1<= level6_c1(30 downto 0) when digit5_c1='1' else level6_c1(62 downto 32);
   digit4_c1<= '1' when level5_c1(30 downto 15) = (15 downto 0 => sozb_c1) else '0';
   level4_c1<= level5_c1(14 downto 0) when digit4_c1='1' else level5_c1(30 downto 16);
   digit3_c2<= '1' when level4_c2(14 downto 7) = (7 downto 0 => sozb_c2) else '0';
   level3_c2<= level4_c2(6 downto 0) when digit3_c2='1' else level4_c2(14 downto 8);
   digit2_c2<= '1' when level3_c2(6 downto 3) = (3 downto 0 => sozb_c2) else '0';
   level2_c2<= level3_c2(2 downto 0) when digit2_c2='1' else level3_c2(6 downto 4);
   -- Finish counting with one LUT
   z_c2 <= level2_c2 when OZB_c2='0' else (not level2_c2);
   with z_c2  select  lowBits_c2 <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits_c2 <= digit6_c2 & digit5_c2 & digit4_c2 & digit3_c2 & digit2_c2 & "";
   O <= outHighBits_c2 & lowBits_c2 ;
end architecture;

--------------------------------------------------------------------------------
--                   LeftShifter34_by_max_34_Freq300_uid13
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X S
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter34_by_max_34_Freq300_uid13 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(33 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(67 downto 0)   );
end entity;

architecture arch of LeftShifter34_by_max_34_Freq300_uid13 is
signal ps_c3, ps_c4 :  std_logic_vector(5 downto 0);
signal level0_c0, level0_c1, level0_c2, level0_c3 :  std_logic_vector(33 downto 0);
signal level1_c3 :  std_logic_vector(34 downto 0);
signal level2_c3 :  std_logic_vector(36 downto 0);
signal level3_c3, level3_c4 :  std_logic_vector(40 downto 0);
signal level4_c4 :  std_logic_vector(48 downto 0);
signal level5_c4 :  std_logic_vector(64 downto 0);
signal level6_c4 :  std_logic_vector(96 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               level0_c1 <= level0_c0;
            end if;
            if ce_2 = '1' then
               level0_c2 <= level0_c1;
            end if;
            if ce_3 = '1' then
               level0_c3 <= level0_c2;
            end if;
            if ce_4 = '1' then
               ps_c4 <= ps_c3;
               level3_c4 <= level3_c3;
            end if;
         end if;
      end process;
   ps_c3<= S;
   level0_c0<= X;
   level1_c3<= level0_c3 & (0 downto 0 => '0') when ps_c3(0)= '1' else     (0 downto 0 => '0') & level0_c3;
   level2_c3<= level1_c3 & (1 downto 0 => '0') when ps_c3(1)= '1' else     (1 downto 0 => '0') & level1_c3;
   level3_c3<= level2_c3 & (3 downto 0 => '0') when ps_c3(2)= '1' else     (3 downto 0 => '0') & level2_c3;
   level4_c4<= level3_c4 & (7 downto 0 => '0') when ps_c4(3)= '1' else     (7 downto 0 => '0') & level3_c4;
   level5_c4<= level4_c4 & (15 downto 0 => '0') when ps_c4(4)= '1' else     (15 downto 0 => '0') & level4_c4;
   level6_c4<= level5_c4 & (31 downto 0 => '0') when ps_c4(5)= '1' else     (31 downto 0 => '0') & level5_c4;
   R <= level6_c4(67 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          InvA0Table_Freq300_uid15
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InvA0Table_Freq300_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of InvA0Table_Freq300_uid15 is
signal Y0_c0 :  std_logic_vector(11 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c0 :  std_logic_vector(11 downto 0);
begin
   with X  select  Y0_c0 <= 
      "100000000000" when "00000000000",
      "100000000000" when "00000000001",
      "011111111111" when "00000000010",
      "011111111110" when "00000000011",
      "011111111101" when "00000000100",
      "011111111100" when "00000000101",
      "011111111011" when "00000000110",
      "011111111010" when "00000000111",
      "011111111001" when "00000001000",
      "011111111000" when "00000001001",
      "011111110111" when "00000001010",
      "011111110110" when "00000001011",
      "011111110101" when "00000001100",
      "011111110100" when "00000001101",
      "011111110011" when "00000001110",
      "011111110010" when "00000001111",
      "011111110001" when "00000010000",
      "011111110000" when "00000010001",
      "011111101111" when "00000010010",
      "011111101110" when "00000010011",
      "011111101101" when "00000010100",
      "011111101100" when "00000010101",
      "011111101011" when "00000010110",
      "011111101010" when "00000010111",
      "011111101001" when "00000011000",
      "011111101000" when "00000011001",
      "011111100111" when "00000011010",
      "011111100110" when "00000011011",
      "011111100101" when "00000011100",
      "011111100100" when "00000011101",
      "011111100011" when "00000011110",
      "011111100010" when "00000011111",
      "011111100001" when "00000100000",
      "011111100000" when "00000100001",
      "011111011111" when "00000100010",
      "011111011110" when "00000100011",
      "011111011101" when "00000100100",
      "011111011100" when "00000100101",
      "011111011011" when "00000100110",
      "011111011010" when "00000100111",
      "011111011001" when "00000101000",
      "011111011000" when "00000101001",
      "011111010111" when "00000101010",
      "011111010110" when "00000101011",
      "011111010101" when "00000101100",
      "011111010100" when "00000101101",
      "011111010100" when "00000101110",
      "011111010011" when "00000101111",
      "011111010010" when "00000110000",
      "011111010001" when "00000110001",
      "011111010000" when "00000110010",
      "011111001111" when "00000110011",
      "011111001110" when "00000110100",
      "011111001101" when "00000110101",
      "011111001100" when "00000110110",
      "011111001011" when "00000110111",
      "011111001010" when "00000111000",
      "011111001001" when "00000111001",
      "011111001000" when "00000111010",
      "011111000111" when "00000111011",
      "011111000110" when "00000111100",
      "011111000101" when "00000111101",
      "011111000100" when "00000111110",
      "011111000011" when "00000111111",
      "011111000010" when "00001000000",
      "011111000001" when "00001000001",
      "011111000001" when "00001000010",
      "011111000000" when "00001000011",
      "011110111111" when "00001000100",
      "011110111110" when "00001000101",
      "011110111101" when "00001000110",
      "011110111100" when "00001000111",
      "011110111011" when "00001001000",
      "011110111010" when "00001001001",
      "011110111001" when "00001001010",
      "011110111000" when "00001001011",
      "011110110111" when "00001001100",
      "011110110110" when "00001001101",
      "011110110101" when "00001001110",
      "011110110100" when "00001001111",
      "011110110100" when "00001010000",
      "011110110011" when "00001010001",
      "011110110010" when "00001010010",
      "011110110001" when "00001010011",
      "011110110000" when "00001010100",
      "011110101111" when "00001010101",
      "011110101110" when "00001010110",
      "011110101101" when "00001010111",
      "011110101100" when "00001011000",
      "011110101011" when "00001011001",
      "011110101010" when "00001011010",
      "011110101001" when "00001011011",
      "011110101000" when "00001011100",
      "011110101000" when "00001011101",
      "011110100111" when "00001011110",
      "011110100110" when "00001011111",
      "011110100101" when "00001100000",
      "011110100100" when "00001100001",
      "011110100011" when "00001100010",
      "011110100010" when "00001100011",
      "011110100001" when "00001100100",
      "011110100000" when "00001100101",
      "011110011111" when "00001100110",
      "011110011110" when "00001100111",
      "011110011110" when "00001101000",
      "011110011101" when "00001101001",
      "011110011100" when "00001101010",
      "011110011011" when "00001101011",
      "011110011010" when "00001101100",
      "011110011001" when "00001101101",
      "011110011000" when "00001101110",
      "011110010111" when "00001101111",
      "011110010110" when "00001110000",
      "011110010101" when "00001110001",
      "011110010101" when "00001110010",
      "011110010100" when "00001110011",
      "011110010011" when "00001110100",
      "011110010010" when "00001110101",
      "011110010001" when "00001110110",
      "011110010000" when "00001110111",
      "011110001111" when "00001111000",
      "011110001110" when "00001111001",
      "011110001101" when "00001111010",
      "011110001100" when "00001111011",
      "011110001100" when "00001111100",
      "011110001011" when "00001111101",
      "011110001010" when "00001111110",
      "011110001001" when "00001111111",
      "011110001000" when "00010000000",
      "011110000111" when "00010000001",
      "011110000110" when "00010000010",
      "011110000101" when "00010000011",
      "011110000100" when "00010000100",
      "011110000100" when "00010000101",
      "011110000011" when "00010000110",
      "011110000010" when "00010000111",
      "011110000001" when "00010001000",
      "011110000000" when "00010001001",
      "011101111111" when "00010001010",
      "011101111110" when "00010001011",
      "011101111101" when "00010001100",
      "011101111101" when "00010001101",
      "011101111100" when "00010001110",
      "011101111011" when "00010001111",
      "011101111010" when "00010010000",
      "011101111001" when "00010010001",
      "011101111000" when "00010010010",
      "011101110111" when "00010010011",
      "011101110110" when "00010010100",
      "011101110110" when "00010010101",
      "011101110101" when "00010010110",
      "011101110100" when "00010010111",
      "011101110011" when "00010011000",
      "011101110010" when "00010011001",
      "011101110001" when "00010011010",
      "011101110000" when "00010011011",
      "011101110000" when "00010011100",
      "011101101111" when "00010011101",
      "011101101110" when "00010011110",
      "011101101101" when "00010011111",
      "011101101100" when "00010100000",
      "011101101011" when "00010100001",
      "011101101010" when "00010100010",
      "011101101010" when "00010100011",
      "011101101001" when "00010100100",
      "011101101000" when "00010100101",
      "011101100111" when "00010100110",
      "011101100110" when "00010100111",
      "011101100101" when "00010101000",
      "011101100100" when "00010101001",
      "011101100100" when "00010101010",
      "011101100011" when "00010101011",
      "011101100010" when "00010101100",
      "011101100001" when "00010101101",
      "011101100000" when "00010101110",
      "011101011111" when "00010101111",
      "011101011110" when "00010110000",
      "011101011110" when "00010110001",
      "011101011101" when "00010110010",
      "011101011100" when "00010110011",
      "011101011011" when "00010110100",
      "011101011010" when "00010110101",
      "011101011001" when "00010110110",
      "011101011001" when "00010110111",
      "011101011000" when "00010111000",
      "011101010111" when "00010111001",
      "011101010110" when "00010111010",
      "011101010101" when "00010111011",
      "011101010100" when "00010111100",
      "011101010011" when "00010111101",
      "011101010011" when "00010111110",
      "011101010010" when "00010111111",
      "011101010001" when "00011000000",
      "011101010000" when "00011000001",
      "011101001111" when "00011000010",
      "011101001110" when "00011000011",
      "011101001110" when "00011000100",
      "011101001101" when "00011000101",
      "011101001100" when "00011000110",
      "011101001011" when "00011000111",
      "011101001010" when "00011001000",
      "011101001001" when "00011001001",
      "011101001001" when "00011001010",
      "011101001000" when "00011001011",
      "011101000111" when "00011001100",
      "011101000110" when "00011001101",
      "011101000101" when "00011001110",
      "011101000101" when "00011001111",
      "011101000100" when "00011010000",
      "011101000011" when "00011010001",
      "011101000010" when "00011010010",
      "011101000001" when "00011010011",
      "011101000000" when "00011010100",
      "011101000000" when "00011010101",
      "011100111111" when "00011010110",
      "011100111110" when "00011010111",
      "011100111101" when "00011011000",
      "011100111100" when "00011011001",
      "011100111011" when "00011011010",
      "011100111011" when "00011011011",
      "011100111010" when "00011011100",
      "011100111001" when "00011011101",
      "011100111000" when "00011011110",
      "011100110111" when "00011011111",
      "011100110111" when "00011100000",
      "011100110110" when "00011100001",
      "011100110101" when "00011100010",
      "011100110100" when "00011100011",
      "011100110011" when "00011100100",
      "011100110011" when "00011100101",
      "011100110010" when "00011100110",
      "011100110001" when "00011100111",
      "011100110000" when "00011101000",
      "011100101111" when "00011101001",
      "011100101110" when "00011101010",
      "011100101110" when "00011101011",
      "011100101101" when "00011101100",
      "011100101100" when "00011101101",
      "011100101011" when "00011101110",
      "011100101010" when "00011101111",
      "011100101010" when "00011110000",
      "011100101001" when "00011110001",
      "011100101000" when "00011110010",
      "011100100111" when "00011110011",
      "011100100110" when "00011110100",
      "011100100110" when "00011110101",
      "011100100101" when "00011110110",
      "011100100100" when "00011110111",
      "011100100011" when "00011111000",
      "011100100010" when "00011111001",
      "011100100010" when "00011111010",
      "011100100001" when "00011111011",
      "011100100000" when "00011111100",
      "011100011111" when "00011111101",
      "011100011111" when "00011111110",
      "011100011110" when "00011111111",
      "011100011101" when "00100000000",
      "011100011100" when "00100000001",
      "011100011011" when "00100000010",
      "011100011011" when "00100000011",
      "011100011010" when "00100000100",
      "011100011001" when "00100000101",
      "011100011000" when "00100000110",
      "011100010111" when "00100000111",
      "011100010111" when "00100001000",
      "011100010110" when "00100001001",
      "011100010101" when "00100001010",
      "011100010100" when "00100001011",
      "011100010100" when "00100001100",
      "011100010011" when "00100001101",
      "011100010010" when "00100001110",
      "011100010001" when "00100001111",
      "011100010000" when "00100010000",
      "011100010000" when "00100010001",
      "011100001111" when "00100010010",
      "011100001110" when "00100010011",
      "011100001101" when "00100010100",
      "011100001101" when "00100010101",
      "011100001100" when "00100010110",
      "011100001011" when "00100010111",
      "011100001010" when "00100011000",
      "011100001001" when "00100011001",
      "011100001001" when "00100011010",
      "011100001000" when "00100011011",
      "011100000111" when "00100011100",
      "011100000110" when "00100011101",
      "011100000110" when "00100011110",
      "011100000101" when "00100011111",
      "011100000100" when "00100100000",
      "011100000011" when "00100100001",
      "011100000010" when "00100100010",
      "011100000010" when "00100100011",
      "011100000001" when "00100100100",
      "011100000000" when "00100100101",
      "011011111111" when "00100100110",
      "011011111111" when "00100100111",
      "011011111110" when "00100101000",
      "011011111101" when "00100101001",
      "011011111100" when "00100101010",
      "011011111100" when "00100101011",
      "011011111011" when "00100101100",
      "011011111010" when "00100101101",
      "011011111001" when "00100101110",
      "011011111001" when "00100101111",
      "011011111000" when "00100110000",
      "011011110111" when "00100110001",
      "011011110110" when "00100110010",
      "011011110110" when "00100110011",
      "011011110101" when "00100110100",
      "011011110100" when "00100110101",
      "011011110011" when "00100110110",
      "011011110011" when "00100110111",
      "011011110010" when "00100111000",
      "011011110001" when "00100111001",
      "011011110000" when "00100111010",
      "011011101111" when "00100111011",
      "011011101111" when "00100111100",
      "011011101110" when "00100111101",
      "011011101101" when "00100111110",
      "011011101100" when "00100111111",
      "011011101100" when "00101000000",
      "011011101011" when "00101000001",
      "011011101010" when "00101000010",
      "011011101010" when "00101000011",
      "011011101001" when "00101000100",
      "011011101000" when "00101000101",
      "011011100111" when "00101000110",
      "011011100111" when "00101000111",
      "011011100110" when "00101001000",
      "011011100101" when "00101001001",
      "011011100100" when "00101001010",
      "011011100100" when "00101001011",
      "011011100011" when "00101001100",
      "011011100010" when "00101001101",
      "011011100001" when "00101001110",
      "011011100001" when "00101001111",
      "011011100000" when "00101010000",
      "011011011111" when "00101010001",
      "011011011110" when "00101010010",
      "011011011110" when "00101010011",
      "011011011101" when "00101010100",
      "011011011100" when "00101010101",
      "011011011011" when "00101010110",
      "011011011011" when "00101010111",
      "011011011010" when "00101011000",
      "011011011001" when "00101011001",
      "011011011001" when "00101011010",
      "011011011000" when "00101011011",
      "011011010111" when "00101011100",
      "011011010110" when "00101011101",
      "011011010110" when "00101011110",
      "011011010101" when "00101011111",
      "011011010100" when "00101100000",
      "011011010011" when "00101100001",
      "011011010011" when "00101100010",
      "011011010010" when "00101100011",
      "011011010001" when "00101100100",
      "011011010000" when "00101100101",
      "011011010000" when "00101100110",
      "011011001111" when "00101100111",
      "011011001110" when "00101101000",
      "011011001110" when "00101101001",
      "011011001101" when "00101101010",
      "011011001100" when "00101101011",
      "011011001011" when "00101101100",
      "011011001011" when "00101101101",
      "011011001010" when "00101101110",
      "011011001001" when "00101101111",
      "011011001001" when "00101110000",
      "011011001000" when "00101110001",
      "011011000111" when "00101110010",
      "011011000110" when "00101110011",
      "011011000110" when "00101110100",
      "011011000101" when "00101110101",
      "011011000100" when "00101110110",
      "011011000100" when "00101110111",
      "011011000011" when "00101111000",
      "011011000010" when "00101111001",
      "011011000001" when "00101111010",
      "011011000001" when "00101111011",
      "011011000000" when "00101111100",
      "011010111111" when "00101111101",
      "011010111111" when "00101111110",
      "011010111110" when "00101111111",
      "011010111101" when "00110000000",
      "011010111100" when "00110000001",
      "011010111100" when "00110000010",
      "011010111011" when "00110000011",
      "011010111010" when "00110000100",
      "011010111010" when "00110000101",
      "011010111001" when "00110000110",
      "011010111000" when "00110000111",
      "011010110111" when "00110001000",
      "011010110111" when "00110001001",
      "011010110110" when "00110001010",
      "011010110101" when "00110001011",
      "011010110101" when "00110001100",
      "011010110100" when "00110001101",
      "011010110011" when "00110001110",
      "011010110011" when "00110001111",
      "011010110010" when "00110010000",
      "011010110001" when "00110010001",
      "011010110000" when "00110010010",
      "011010110000" when "00110010011",
      "011010101111" when "00110010100",
      "011010101110" when "00110010101",
      "011010101110" when "00110010110",
      "011010101101" when "00110010111",
      "011010101100" when "00110011000",
      "011010101100" when "00110011001",
      "011010101011" when "00110011010",
      "011010101010" when "00110011011",
      "011010101010" when "00110011100",
      "011010101001" when "00110011101",
      "011010101000" when "00110011110",
      "011010100111" when "00110011111",
      "011010100111" when "00110100000",
      "011010100110" when "00110100001",
      "011010100101" when "00110100010",
      "011010100101" when "00110100011",
      "011010100100" when "00110100100",
      "011010100011" when "00110100101",
      "011010100011" when "00110100110",
      "011010100010" when "00110100111",
      "011010100001" when "00110101000",
      "011010100001" when "00110101001",
      "011010100000" when "00110101010",
      "011010011111" when "00110101011",
      "011010011110" when "00110101100",
      "011010011110" when "00110101101",
      "011010011101" when "00110101110",
      "011010011100" when "00110101111",
      "011010011100" when "00110110000",
      "011010011011" when "00110110001",
      "011010011010" when "00110110010",
      "011010011010" when "00110110011",
      "011010011001" when "00110110100",
      "011010011000" when "00110110101",
      "011010011000" when "00110110110",
      "011010010111" when "00110110111",
      "011010010110" when "00110111000",
      "011010010110" when "00110111001",
      "011010010101" when "00110111010",
      "011010010100" when "00110111011",
      "011010010100" when "00110111100",
      "011010010011" when "00110111101",
      "011010010010" when "00110111110",
      "011010010010" when "00110111111",
      "011010010001" when "00111000000",
      "011010010000" when "00111000001",
      "011010010000" when "00111000010",
      "011010001111" when "00111000011",
      "011010001110" when "00111000100",
      "011010001110" when "00111000101",
      "011010001101" when "00111000110",
      "011010001100" when "00111000111",
      "011010001100" when "00111001000",
      "011010001011" when "00111001001",
      "011010001010" when "00111001010",
      "011010001010" when "00111001011",
      "011010001001" when "00111001100",
      "011010001000" when "00111001101",
      "011010001000" when "00111001110",
      "011010000111" when "00111001111",
      "011010000110" when "00111010000",
      "011010000110" when "00111010001",
      "011010000101" when "00111010010",
      "011010000100" when "00111010011",
      "011010000100" when "00111010100",
      "011010000011" when "00111010101",
      "011010000010" when "00111010110",
      "011010000010" when "00111010111",
      "011010000001" when "00111011000",
      "011010000000" when "00111011001",
      "011010000000" when "00111011010",
      "011001111111" when "00111011011",
      "011001111110" when "00111011100",
      "011001111110" when "00111011101",
      "011001111101" when "00111011110",
      "011001111100" when "00111011111",
      "011001111100" when "00111100000",
      "011001111011" when "00111100001",
      "011001111010" when "00111100010",
      "011001111010" when "00111100011",
      "011001111001" when "00111100100",
      "011001111000" when "00111100101",
      "011001111000" when "00111100110",
      "011001110111" when "00111100111",
      "011001110110" when "00111101000",
      "011001110110" when "00111101001",
      "011001110101" when "00111101010",
      "011001110100" when "00111101011",
      "011001110100" when "00111101100",
      "011001110011" when "00111101101",
      "011001110011" when "00111101110",
      "011001110010" when "00111101111",
      "011001110001" when "00111110000",
      "011001110001" when "00111110001",
      "011001110000" when "00111110010",
      "011001101111" when "00111110011",
      "011001101111" when "00111110100",
      "011001101110" when "00111110101",
      "011001101101" when "00111110110",
      "011001101101" when "00111110111",
      "011001101100" when "00111111000",
      "011001101011" when "00111111001",
      "011001101011" when "00111111010",
      "011001101010" when "00111111011",
      "011001101001" when "00111111100",
      "011001101001" when "00111111101",
      "011001101000" when "00111111110",
      "011001101000" when "00111111111",
      "011001100111" when "01000000000",
      "011001100110" when "01000000001",
      "011001100110" when "01000000010",
      "011001100101" when "01000000011",
      "011001100100" when "01000000100",
      "011001100100" when "01000000101",
      "011001100011" when "01000000110",
      "011001100010" when "01000000111",
      "011001100010" when "01000001000",
      "011001100001" when "01000001001",
      "011001100001" when "01000001010",
      "011001100000" when "01000001011",
      "011001011111" when "01000001100",
      "011001011111" when "01000001101",
      "011001011110" when "01000001110",
      "011001011101" when "01000001111",
      "011001011101" when "01000010000",
      "011001011100" when "01000010001",
      "011001011011" when "01000010010",
      "011001011011" when "01000010011",
      "011001011010" when "01000010100",
      "011001011010" when "01000010101",
      "011001011001" when "01000010110",
      "011001011000" when "01000010111",
      "011001011000" when "01000011000",
      "011001010111" when "01000011001",
      "011001010110" when "01000011010",
      "011001010110" when "01000011011",
      "011001010101" when "01000011100",
      "011001010101" when "01000011101",
      "011001010100" when "01000011110",
      "011001010011" when "01000011111",
      "011001010011" when "01000100000",
      "011001010010" when "01000100001",
      "011001010001" when "01000100010",
      "011001010001" when "01000100011",
      "011001010000" when "01000100100",
      "011001010000" when "01000100101",
      "011001001111" when "01000100110",
      "011001001110" when "01000100111",
      "011001001110" when "01000101000",
      "011001001101" when "01000101001",
      "011001001100" when "01000101010",
      "011001001100" when "01000101011",
      "011001001011" when "01000101100",
      "011001001011" when "01000101101",
      "011001001010" when "01000101110",
      "011001001001" when "01000101111",
      "011001001001" when "01000110000",
      "011001001000" when "01000110001",
      "011001001000" when "01000110010",
      "011001000111" when "01000110011",
      "011001000110" when "01000110100",
      "011001000110" when "01000110101",
      "011001000101" when "01000110110",
      "011001000100" when "01000110111",
      "011001000100" when "01000111000",
      "011001000011" when "01000111001",
      "011001000011" when "01000111010",
      "011001000010" when "01000111011",
      "011001000001" when "01000111100",
      "011001000001" when "01000111101",
      "011001000000" when "01000111110",
      "011001000000" when "01000111111",
      "011000111111" when "01001000000",
      "011000111110" when "01001000001",
      "011000111110" when "01001000010",
      "011000111101" when "01001000011",
      "011000111101" when "01001000100",
      "011000111100" when "01001000101",
      "011000111011" when "01001000110",
      "011000111011" when "01001000111",
      "011000111010" when "01001001000",
      "011000111001" when "01001001001",
      "011000111001" when "01001001010",
      "011000111000" when "01001001011",
      "011000111000" when "01001001100",
      "011000110111" when "01001001101",
      "011000110110" when "01001001110",
      "011000110110" when "01001001111",
      "011000110101" when "01001010000",
      "011000110101" when "01001010001",
      "011000110100" when "01001010010",
      "011000110011" when "01001010011",
      "011000110011" when "01001010100",
      "011000110010" when "01001010101",
      "011000110010" when "01001010110",
      "011000110001" when "01001010111",
      "011000110000" when "01001011000",
      "011000110000" when "01001011001",
      "011000101111" when "01001011010",
      "011000101111" when "01001011011",
      "011000101110" when "01001011100",
      "011000101101" when "01001011101",
      "011000101101" when "01001011110",
      "011000101100" when "01001011111",
      "011000101100" when "01001100000",
      "011000101011" when "01001100001",
      "011000101010" when "01001100010",
      "011000101010" when "01001100011",
      "011000101001" when "01001100100",
      "011000101001" when "01001100101",
      "011000101000" when "01001100110",
      "011000101000" when "01001100111",
      "011000100111" when "01001101000",
      "011000100110" when "01001101001",
      "011000100110" when "01001101010",
      "011000100101" when "01001101011",
      "011000100101" when "01001101100",
      "011000100100" when "01001101101",
      "011000100011" when "01001101110",
      "011000100011" when "01001101111",
      "011000100010" when "01001110000",
      "011000100010" when "01001110001",
      "011000100001" when "01001110010",
      "011000100000" when "01001110011",
      "011000100000" when "01001110100",
      "011000011111" when "01001110101",
      "011000011111" when "01001110110",
      "011000011110" when "01001110111",
      "011000011110" when "01001111000",
      "011000011101" when "01001111001",
      "011000011100" when "01001111010",
      "011000011100" when "01001111011",
      "011000011011" when "01001111100",
      "011000011011" when "01001111101",
      "011000011010" when "01001111110",
      "011000011001" when "01001111111",
      "011000011001" when "01010000000",
      "011000011000" when "01010000001",
      "011000011000" when "01010000010",
      "011000010111" when "01010000011",
      "011000010111" when "01010000100",
      "011000010110" when "01010000101",
      "011000010101" when "01010000110",
      "011000010101" when "01010000111",
      "011000010100" when "01010001000",
      "011000010100" when "01010001001",
      "011000010011" when "01010001010",
      "011000010011" when "01010001011",
      "011000010010" when "01010001100",
      "011000010001" when "01010001101",
      "011000010001" when "01010001110",
      "011000010000" when "01010001111",
      "011000010000" when "01010010000",
      "011000001111" when "01010010001",
      "011000001111" when "01010010010",
      "011000001110" when "01010010011",
      "011000001101" when "01010010100",
      "011000001101" when "01010010101",
      "011000001100" when "01010010110",
      "011000001100" when "01010010111",
      "011000001011" when "01010011000",
      "011000001011" when "01010011001",
      "011000001010" when "01010011010",
      "011000001001" when "01010011011",
      "011000001001" when "01010011100",
      "011000001000" when "01010011101",
      "011000001000" when "01010011110",
      "011000000111" when "01010011111",
      "011000000111" when "01010100000",
      "011000000110" when "01010100001",
      "011000000101" when "01010100010",
      "011000000101" when "01010100011",
      "011000000100" when "01010100100",
      "011000000100" when "01010100101",
      "011000000011" when "01010100110",
      "011000000011" when "01010100111",
      "011000000010" when "01010101000",
      "011000000001" when "01010101001",
      "011000000001" when "01010101010",
      "011000000000" when "01010101011",
      "011000000000" when "01010101100",
      "010111111111" when "01010101101",
      "010111111111" when "01010101110",
      "010111111110" when "01010101111",
      "010111111110" when "01010110000",
      "010111111101" when "01010110001",
      "010111111100" when "01010110010",
      "010111111100" when "01010110011",
      "010111111011" when "01010110100",
      "010111111011" when "01010110101",
      "010111111010" when "01010110110",
      "010111111010" when "01010110111",
      "010111111001" when "01010111000",
      "010111111000" when "01010111001",
      "010111111000" when "01010111010",
      "010111110111" when "01010111011",
      "010111110111" when "01010111100",
      "010111110110" when "01010111101",
      "010111110110" when "01010111110",
      "010111110101" when "01010111111",
      "010111110101" when "01011000000",
      "010111110100" when "01011000001",
      "010111110011" when "01011000010",
      "010111110011" when "01011000011",
      "010111110010" when "01011000100",
      "010111110010" when "01011000101",
      "010111110001" when "01011000110",
      "010111110001" when "01011000111",
      "010111110000" when "01011001000",
      "010111110000" when "01011001001",
      "010111101111" when "01011001010",
      "010111101111" when "01011001011",
      "010111101110" when "01011001100",
      "010111101101" when "01011001101",
      "010111101101" when "01011001110",
      "010111101100" when "01011001111",
      "010111101100" when "01011010000",
      "010111101011" when "01011010001",
      "010111101011" when "01011010010",
      "010111101010" when "01011010011",
      "010111101010" when "01011010100",
      "010111101001" when "01011010101",
      "010111101001" when "01011010110",
      "010111101000" when "01011010111",
      "010111100111" when "01011011000",
      "010111100111" when "01011011001",
      "010111100110" when "01011011010",
      "010111100110" when "01011011011",
      "010111100101" when "01011011100",
      "010111100101" when "01011011101",
      "010111100100" when "01011011110",
      "010111100100" when "01011011111",
      "010111100011" when "01011100000",
      "010111100011" when "01011100001",
      "010111100010" when "01011100010",
      "010111100001" when "01011100011",
      "010111100001" when "01011100100",
      "010111100000" when "01011100101",
      "010111100000" when "01011100110",
      "010111011111" when "01011100111",
      "010111011111" when "01011101000",
      "010111011110" when "01011101001",
      "010111011110" when "01011101010",
      "010111011101" when "01011101011",
      "010111011101" when "01011101100",
      "010111011100" when "01011101101",
      "010111011100" when "01011101110",
      "010111011011" when "01011101111",
      "010111011010" when "01011110000",
      "010111011010" when "01011110001",
      "010111011001" when "01011110010",
      "010111011001" when "01011110011",
      "010111011000" when "01011110100",
      "010111011000" when "01011110101",
      "010111010111" when "01011110110",
      "010111010111" when "01011110111",
      "010111010110" when "01011111000",
      "010111010110" when "01011111001",
      "010111010101" when "01011111010",
      "010111010101" when "01011111011",
      "010111010100" when "01011111100",
      "010111010100" when "01011111101",
      "010111010011" when "01011111110",
      "010111010010" when "01011111111",
      "010111010010" when "01100000000",
      "010111010001" when "01100000001",
      "010111010001" when "01100000010",
      "010111010000" when "01100000011",
      "010111010000" when "01100000100",
      "010111001111" when "01100000101",
      "010111001111" when "01100000110",
      "010111001110" when "01100000111",
      "010111001110" when "01100001000",
      "010111001101" when "01100001001",
      "010111001101" when "01100001010",
      "010111001100" when "01100001011",
      "010111001100" when "01100001100",
      "010111001011" when "01100001101",
      "010111001011" when "01100001110",
      "010111001010" when "01100001111",
      "010111001010" when "01100010000",
      "010111001001" when "01100010001",
      "010111001000" when "01100010010",
      "010111001000" when "01100010011",
      "010111000111" when "01100010100",
      "010111000111" when "01100010101",
      "010111000110" when "01100010110",
      "010111000110" when "01100010111",
      "010111000101" when "01100011000",
      "010111000101" when "01100011001",
      "010111000100" when "01100011010",
      "010111000100" when "01100011011",
      "010111000011" when "01100011100",
      "010111000011" when "01100011101",
      "010111000010" when "01100011110",
      "010111000010" when "01100011111",
      "010111000001" when "01100100000",
      "010111000001" when "01100100001",
      "010111000000" when "01100100010",
      "010111000000" when "01100100011",
      "010110111111" when "01100100100",
      "010110111111" when "01100100101",
      "010110111110" when "01100100110",
      "010110111110" when "01100100111",
      "010110111101" when "01100101000",
      "010110111101" when "01100101001",
      "010110111100" when "01100101010",
      "010110111100" when "01100101011",
      "010110111011" when "01100101100",
      "010110111011" when "01100101101",
      "010110111010" when "01100101110",
      "010110111010" when "01100101111",
      "010110111001" when "01100110000",
      "010110111000" when "01100110001",
      "010110111000" when "01100110010",
      "010110110111" when "01100110011",
      "010110110111" when "01100110100",
      "010110110110" when "01100110101",
      "010110110110" when "01100110110",
      "010110110101" when "01100110111",
      "010110110101" when "01100111000",
      "010110110100" when "01100111001",
      "010110110100" when "01100111010",
      "010110110011" when "01100111011",
      "010110110011" when "01100111100",
      "010110110010" when "01100111101",
      "010110110010" when "01100111110",
      "010110110001" when "01100111111",
      "010110110001" when "01101000000",
      "010110110000" when "01101000001",
      "010110110000" when "01101000010",
      "010110101111" when "01101000011",
      "010110101111" when "01101000100",
      "010110101110" when "01101000101",
      "010110101110" when "01101000110",
      "010110101101" when "01101000111",
      "010110101101" when "01101001000",
      "010110101100" when "01101001001",
      "010110101100" when "01101001010",
      "010110101011" when "01101001011",
      "010110101011" when "01101001100",
      "010110101010" when "01101001101",
      "010110101010" when "01101001110",
      "010110101001" when "01101001111",
      "010110101001" when "01101010000",
      "010110101000" when "01101010001",
      "010110101000" when "01101010010",
      "010110100111" when "01101010011",
      "010110100111" when "01101010100",
      "010110100110" when "01101010101",
      "010110100110" when "01101010110",
      "010110100101" when "01101010111",
      "010110100101" when "01101011000",
      "010110100100" when "01101011001",
      "010110100100" when "01101011010",
      "010110100011" when "01101011011",
      "010110100011" when "01101011100",
      "010110100010" when "01101011101",
      "010110100010" when "01101011110",
      "010110100001" when "01101011111",
      "010110100001" when "01101100000",
      "010110100000" when "01101100001",
      "010110100000" when "01101100010",
      "010110011111" when "01101100011",
      "010110011111" when "01101100100",
      "010110011110" when "01101100101",
      "010110011110" when "01101100110",
      "010110011101" when "01101100111",
      "010110011101" when "01101101000",
      "010110011100" when "01101101001",
      "010110011100" when "01101101010",
      "010110011011" when "01101101011",
      "010110011011" when "01101101100",
      "010110011010" when "01101101101",
      "010110011010" when "01101101110",
      "010110011001" when "01101101111",
      "010110011001" when "01101110000",
      "010110011000" when "01101110001",
      "010110011000" when "01101110010",
      "010110011000" when "01101110011",
      "010110010111" when "01101110100",
      "010110010111" when "01101110101",
      "010110010110" when "01101110110",
      "010110010110" when "01101110111",
      "010110010101" when "01101111000",
      "010110010101" when "01101111001",
      "010110010100" when "01101111010",
      "010110010100" when "01101111011",
      "010110010011" when "01101111100",
      "010110010011" when "01101111101",
      "010110010010" when "01101111110",
      "010110010010" when "01101111111",
      "010110010001" when "01110000000",
      "010110010001" when "01110000001",
      "010110010000" when "01110000010",
      "010110010000" when "01110000011",
      "010110001111" when "01110000100",
      "010110001111" when "01110000101",
      "010110001110" when "01110000110",
      "010110001110" when "01110000111",
      "010110001101" when "01110001000",
      "010110001101" when "01110001001",
      "010110001100" when "01110001010",
      "010110001100" when "01110001011",
      "010110001011" when "01110001100",
      "010110001011" when "01110001101",
      "010110001010" when "01110001110",
      "010110001010" when "01110001111",
      "010110001001" when "01110010000",
      "010110001001" when "01110010001",
      "010110001001" when "01110010010",
      "010110001000" when "01110010011",
      "010110001000" when "01110010100",
      "010110000111" when "01110010101",
      "010110000111" when "01110010110",
      "010110000110" when "01110010111",
      "010110000110" when "01110011000",
      "010110000101" when "01110011001",
      "010110000101" when "01110011010",
      "010110000100" when "01110011011",
      "010110000100" when "01110011100",
      "010110000011" when "01110011101",
      "010110000011" when "01110011110",
      "010110000010" when "01110011111",
      "010110000010" when "01110100000",
      "010110000001" when "01110100001",
      "010110000001" when "01110100010",
      "010110000000" when "01110100011",
      "010110000000" when "01110100100",
      "010110000000" when "01110100101",
      "010101111111" when "01110100110",
      "010101111111" when "01110100111",
      "010101111110" when "01110101000",
      "010101111110" when "01110101001",
      "010101111101" when "01110101010",
      "010101111101" when "01110101011",
      "010101111100" when "01110101100",
      "010101111100" when "01110101101",
      "010101111011" when "01110101110",
      "010101111011" when "01110101111",
      "010101111010" when "01110110000",
      "010101111010" when "01110110001",
      "010101111001" when "01110110010",
      "010101111001" when "01110110011",
      "010101111000" when "01110110100",
      "010101111000" when "01110110101",
      "010101111000" when "01110110110",
      "010101110111" when "01110110111",
      "010101110111" when "01110111000",
      "010101110110" when "01110111001",
      "010101110110" when "01110111010",
      "010101110101" when "01110111011",
      "010101110101" when "01110111100",
      "010101110100" when "01110111101",
      "010101110100" when "01110111110",
      "010101110011" when "01110111111",
      "010101110011" when "01111000000",
      "010101110010" when "01111000001",
      "010101110010" when "01111000010",
      "010101110001" when "01111000011",
      "010101110001" when "01111000100",
      "010101110001" when "01111000101",
      "010101110000" when "01111000110",
      "010101110000" when "01111000111",
      "010101101111" when "01111001000",
      "010101101111" when "01111001001",
      "010101101110" when "01111001010",
      "010101101110" when "01111001011",
      "010101101101" when "01111001100",
      "010101101101" when "01111001101",
      "010101101100" when "01111001110",
      "010101101100" when "01111001111",
      "010101101100" when "01111010000",
      "010101101011" when "01111010001",
      "010101101011" when "01111010010",
      "010101101010" when "01111010011",
      "010101101010" when "01111010100",
      "010101101001" when "01111010101",
      "010101101001" when "01111010110",
      "010101101000" when "01111010111",
      "010101101000" when "01111011000",
      "010101100111" when "01111011001",
      "010101100111" when "01111011010",
      "010101100110" when "01111011011",
      "010101100110" when "01111011100",
      "010101100110" when "01111011101",
      "010101100101" when "01111011110",
      "010101100101" when "01111011111",
      "010101100100" when "01111100000",
      "010101100100" when "01111100001",
      "010101100011" when "01111100010",
      "010101100011" when "01111100011",
      "010101100010" when "01111100100",
      "010101100010" when "01111100101",
      "010101100001" when "01111100110",
      "010101100001" when "01111100111",
      "010101100001" when "01111101000",
      "010101100000" when "01111101001",
      "010101100000" when "01111101010",
      "010101011111" when "01111101011",
      "010101011111" when "01111101100",
      "010101011110" when "01111101101",
      "010101011110" when "01111101110",
      "010101011101" when "01111101111",
      "010101011101" when "01111110000",
      "010101011101" when "01111110001",
      "010101011100" when "01111110010",
      "010101011100" when "01111110011",
      "010101011011" when "01111110100",
      "010101011011" when "01111110101",
      "010101011010" when "01111110110",
      "010101011010" when "01111110111",
      "010101011001" when "01111111000",
      "010101011001" when "01111111001",
      "010101011001" when "01111111010",
      "010101011000" when "01111111011",
      "010101011000" when "01111111100",
      "010101010111" when "01111111101",
      "010101010111" when "01111111110",
      "010101010110" when "01111111111",
      "101010101011" when "10000000000",
      "101010101010" when "10000000001",
      "101010101001" when "10000000010",
      "101010101001" when "10000000011",
      "101010101000" when "10000000100",
      "101010100111" when "10000000101",
      "101010100110" when "10000000110",
      "101010100101" when "10000000111",
      "101010100100" when "10000001000",
      "101010100011" when "10000001001",
      "101010100010" when "10000001010",
      "101010100001" when "10000001011",
      "101010100001" when "10000001100",
      "101010100000" when "10000001101",
      "101010011111" when "10000001110",
      "101010011110" when "10000001111",
      "101010011101" when "10000010000",
      "101010011100" when "10000010001",
      "101010011011" when "10000010010",
      "101010011010" when "10000010011",
      "101010011010" when "10000010100",
      "101010011001" when "10000010101",
      "101010011000" when "10000010110",
      "101010010111" when "10000010111",
      "101010010110" when "10000011000",
      "101010010101" when "10000011001",
      "101010010100" when "10000011010",
      "101010010011" when "10000011011",
      "101010010011" when "10000011100",
      "101010010010" when "10000011101",
      "101010010001" when "10000011110",
      "101010010000" when "10000011111",
      "101010001111" when "10000100000",
      "101010001110" when "10000100001",
      "101010001101" when "10000100010",
      "101010001100" when "10000100011",
      "101010001100" when "10000100100",
      "101010001011" when "10000100101",
      "101010001010" when "10000100110",
      "101010001001" when "10000100111",
      "101010001000" when "10000101000",
      "101010000111" when "10000101001",
      "101010000110" when "10000101010",
      "101010000101" when "10000101011",
      "101010000101" when "10000101100",
      "101010000100" when "10000101101",
      "101010000011" when "10000101110",
      "101010000010" when "10000101111",
      "101010000001" when "10000110000",
      "101010000000" when "10000110001",
      "101001111111" when "10000110010",
      "101001111111" when "10000110011",
      "101001111110" when "10000110100",
      "101001111101" when "10000110101",
      "101001111100" when "10000110110",
      "101001111011" when "10000110111",
      "101001111010" when "10000111000",
      "101001111001" when "10000111001",
      "101001111001" when "10000111010",
      "101001111000" when "10000111011",
      "101001110111" when "10000111100",
      "101001110110" when "10000111101",
      "101001110101" when "10000111110",
      "101001110100" when "10000111111",
      "101001110011" when "10001000000",
      "101001110011" when "10001000001",
      "101001110010" when "10001000010",
      "101001110001" when "10001000011",
      "101001110000" when "10001000100",
      "101001101111" when "10001000101",
      "101001101110" when "10001000110",
      "101001101101" when "10001000111",
      "101001101101" when "10001001000",
      "101001101100" when "10001001001",
      "101001101011" when "10001001010",
      "101001101010" when "10001001011",
      "101001101001" when "10001001100",
      "101001101000" when "10001001101",
      "101001101000" when "10001001110",
      "101001100111" when "10001001111",
      "101001100110" when "10001010000",
      "101001100101" when "10001010001",
      "101001100100" when "10001010010",
      "101001100011" when "10001010011",
      "101001100010" when "10001010100",
      "101001100010" when "10001010101",
      "101001100001" when "10001010110",
      "101001100000" when "10001010111",
      "101001011111" when "10001011000",
      "101001011110" when "10001011001",
      "101001011101" when "10001011010",
      "101001011101" when "10001011011",
      "101001011100" when "10001011100",
      "101001011011" when "10001011101",
      "101001011010" when "10001011110",
      "101001011001" when "10001011111",
      "101001011000" when "10001100000",
      "101001011000" when "10001100001",
      "101001010111" when "10001100010",
      "101001010110" when "10001100011",
      "101001010101" when "10001100100",
      "101001010100" when "10001100101",
      "101001010011" when "10001100110",
      "101001010011" when "10001100111",
      "101001010010" when "10001101000",
      "101001010001" when "10001101001",
      "101001010000" when "10001101010",
      "101001001111" when "10001101011",
      "101001001110" when "10001101100",
      "101001001110" when "10001101101",
      "101001001101" when "10001101110",
      "101001001100" when "10001101111",
      "101001001011" when "10001110000",
      "101001001010" when "10001110001",
      "101001001001" when "10001110010",
      "101001001001" when "10001110011",
      "101001001000" when "10001110100",
      "101001000111" when "10001110101",
      "101001000110" when "10001110110",
      "101001000101" when "10001110111",
      "101001000101" when "10001111000",
      "101001000100" when "10001111001",
      "101001000011" when "10001111010",
      "101001000010" when "10001111011",
      "101001000001" when "10001111100",
      "101001000000" when "10001111101",
      "101001000000" when "10001111110",
      "101000111111" when "10001111111",
      "101000111110" when "10010000000",
      "101000111101" when "10010000001",
      "101000111100" when "10010000010",
      "101000111011" when "10010000011",
      "101000111011" when "10010000100",
      "101000111010" when "10010000101",
      "101000111001" when "10010000110",
      "101000111000" when "10010000111",
      "101000110111" when "10010001000",
      "101000110111" when "10010001001",
      "101000110110" when "10010001010",
      "101000110101" when "10010001011",
      "101000110100" when "10010001100",
      "101000110011" when "10010001101",
      "101000110011" when "10010001110",
      "101000110010" when "10010001111",
      "101000110001" when "10010010000",
      "101000110000" when "10010010001",
      "101000101111" when "10010010010",
      "101000101110" when "10010010011",
      "101000101110" when "10010010100",
      "101000101101" when "10010010101",
      "101000101100" when "10010010110",
      "101000101011" when "10010010111",
      "101000101010" when "10010011000",
      "101000101010" when "10010011001",
      "101000101001" when "10010011010",
      "101000101000" when "10010011011",
      "101000100111" when "10010011100",
      "101000100110" when "10010011101",
      "101000100110" when "10010011110",
      "101000100101" when "10010011111",
      "101000100100" when "10010100000",
      "101000100011" when "10010100001",
      "101000100010" when "10010100010",
      "101000100010" when "10010100011",
      "101000100001" when "10010100100",
      "101000100000" when "10010100101",
      "101000011111" when "10010100110",
      "101000011110" when "10010100111",
      "101000011110" when "10010101000",
      "101000011101" when "10010101001",
      "101000011100" when "10010101010",
      "101000011011" when "10010101011",
      "101000011010" when "10010101100",
      "101000011010" when "10010101101",
      "101000011001" when "10010101110",
      "101000011000" when "10010101111",
      "101000010111" when "10010110000",
      "101000010110" when "10010110001",
      "101000010110" when "10010110010",
      "101000010101" when "10010110011",
      "101000010100" when "10010110100",
      "101000010011" when "10010110101",
      "101000010010" when "10010110110",
      "101000010010" when "10010110111",
      "101000010001" when "10010111000",
      "101000010000" when "10010111001",
      "101000001111" when "10010111010",
      "101000001110" when "10010111011",
      "101000001110" when "10010111100",
      "101000001101" when "10010111101",
      "101000001100" when "10010111110",
      "101000001011" when "10010111111",
      "101000001011" when "10011000000",
      "101000001010" when "10011000001",
      "101000001001" when "10011000010",
      "101000001000" when "10011000011",
      "101000000111" when "10011000100",
      "101000000111" when "10011000101",
      "101000000110" when "10011000110",
      "101000000101" when "10011000111",
      "101000000100" when "10011001000",
      "101000000011" when "10011001001",
      "101000000011" when "10011001010",
      "101000000010" when "10011001011",
      "101000000001" when "10011001100",
      "101000000000" when "10011001101",
      "101000000000" when "10011001110",
      "100111111111" when "10011001111",
      "100111111110" when "10011010000",
      "100111111101" when "10011010001",
      "100111111100" when "10011010010",
      "100111111100" when "10011010011",
      "100111111011" when "10011010100",
      "100111111010" when "10011010101",
      "100111111001" when "10011010110",
      "100111111001" when "10011010111",
      "100111111000" when "10011011000",
      "100111110111" when "10011011001",
      "100111110110" when "10011011010",
      "100111110101" when "10011011011",
      "100111110101" when "10011011100",
      "100111110100" when "10011011101",
      "100111110011" when "10011011110",
      "100111110010" when "10011011111",
      "100111110010" when "10011100000",
      "100111110001" when "10011100001",
      "100111110000" when "10011100010",
      "100111101111" when "10011100011",
      "100111101111" when "10011100100",
      "100111101110" when "10011100101",
      "100111101101" when "10011100110",
      "100111101100" when "10011100111",
      "100111101011" when "10011101000",
      "100111101011" when "10011101001",
      "100111101010" when "10011101010",
      "100111101001" when "10011101011",
      "100111101000" when "10011101100",
      "100111101000" when "10011101101",
      "100111100111" when "10011101110",
      "100111100110" when "10011101111",
      "100111100101" when "10011110000",
      "100111100101" when "10011110001",
      "100111100100" when "10011110010",
      "100111100011" when "10011110011",
      "100111100010" when "10011110100",
      "100111100001" when "10011110101",
      "100111100001" when "10011110110",
      "100111100000" when "10011110111",
      "100111011111" when "10011111000",
      "100111011110" when "10011111001",
      "100111011110" when "10011111010",
      "100111011101" when "10011111011",
      "100111011100" when "10011111100",
      "100111011011" when "10011111101",
      "100111011011" when "10011111110",
      "100111011010" when "10011111111",
      "100111011001" when "10100000000",
      "100111011000" when "10100000001",
      "100111011000" when "10100000010",
      "100111010111" when "10100000011",
      "100111010110" when "10100000100",
      "100111010101" when "10100000101",
      "100111010101" when "10100000110",
      "100111010100" when "10100000111",
      "100111010011" when "10100001000",
      "100111010010" when "10100001001",
      "100111010010" when "10100001010",
      "100111010001" when "10100001011",
      "100111010000" when "10100001100",
      "100111001111" when "10100001101",
      "100111001111" when "10100001110",
      "100111001110" when "10100001111",
      "100111001101" when "10100010000",
      "100111001100" when "10100010001",
      "100111001100" when "10100010010",
      "100111001011" when "10100010011",
      "100111001010" when "10100010100",
      "100111001001" when "10100010101",
      "100111001001" when "10100010110",
      "100111001000" when "10100010111",
      "100111000111" when "10100011000",
      "100111000110" when "10100011001",
      "100111000110" when "10100011010",
      "100111000101" when "10100011011",
      "100111000100" when "10100011100",
      "100111000011" when "10100011101",
      "100111000011" when "10100011110",
      "100111000010" when "10100011111",
      "100111000001" when "10100100000",
      "100111000000" when "10100100001",
      "100111000000" when "10100100010",
      "100110111111" when "10100100011",
      "100110111110" when "10100100100",
      "100110111101" when "10100100101",
      "100110111101" when "10100100110",
      "100110111100" when "10100100111",
      "100110111011" when "10100101000",
      "100110111010" when "10100101001",
      "100110111010" when "10100101010",
      "100110111001" when "10100101011",
      "100110111000" when "10100101100",
      "100110110111" when "10100101101",
      "100110110111" when "10100101110",
      "100110110110" when "10100101111",
      "100110110101" when "10100110000",
      "100110110101" when "10100110001",
      "100110110100" when "10100110010",
      "100110110011" when "10100110011",
      "100110110010" when "10100110100",
      "100110110010" when "10100110101",
      "100110110001" when "10100110110",
      "100110110000" when "10100110111",
      "100110101111" when "10100111000",
      "100110101111" when "10100111001",
      "100110101110" when "10100111010",
      "100110101101" when "10100111011",
      "100110101100" when "10100111100",
      "100110101100" when "10100111101",
      "100110101011" when "10100111110",
      "100110101010" when "10100111111",
      "100110101010" when "10101000000",
      "100110101001" when "10101000001",
      "100110101000" when "10101000010",
      "100110100111" when "10101000011",
      "100110100111" when "10101000100",
      "100110100110" when "10101000101",
      "100110100101" when "10101000110",
      "100110100100" when "10101000111",
      "100110100100" when "10101001000",
      "100110100011" when "10101001001",
      "100110100010" when "10101001010",
      "100110100010" when "10101001011",
      "100110100001" when "10101001100",
      "100110100000" when "10101001101",
      "100110011111" when "10101001110",
      "100110011111" when "10101001111",
      "100110011110" when "10101010000",
      "100110011101" when "10101010001",
      "100110011101" when "10101010010",
      "100110011100" when "10101010011",
      "100110011011" when "10101010100",
      "100110011010" when "10101010101",
      "100110011010" when "10101010110",
      "100110011001" when "10101010111",
      "100110011000" when "10101011000",
      "100110010111" when "10101011001",
      "100110010111" when "10101011010",
      "100110010110" when "10101011011",
      "100110010101" when "10101011100",
      "100110010101" when "10101011101",
      "100110010100" when "10101011110",
      "100110010011" when "10101011111",
      "100110010010" when "10101100000",
      "100110010010" when "10101100001",
      "100110010001" when "10101100010",
      "100110010000" when "10101100011",
      "100110010000" when "10101100100",
      "100110001111" when "10101100101",
      "100110001110" when "10101100110",
      "100110001101" when "10101100111",
      "100110001101" when "10101101000",
      "100110001100" when "10101101001",
      "100110001011" when "10101101010",
      "100110001011" when "10101101011",
      "100110001010" when "10101101100",
      "100110001001" when "10101101101",
      "100110001000" when "10101101110",
      "100110001000" when "10101101111",
      "100110000111" when "10101110000",
      "100110000110" when "10101110001",
      "100110000110" when "10101110010",
      "100110000101" when "10101110011",
      "100110000100" when "10101110100",
      "100110000100" when "10101110101",
      "100110000011" when "10101110110",
      "100110000010" when "10101110111",
      "100110000001" when "10101111000",
      "100110000001" when "10101111001",
      "100110000000" when "10101111010",
      "100101111111" when "10101111011",
      "100101111111" when "10101111100",
      "100101111110" when "10101111101",
      "100101111101" when "10101111110",
      "100101111100" when "10101111111",
      "100101111100" when "10110000000",
      "100101111011" when "10110000001",
      "100101111010" when "10110000010",
      "100101111010" when "10110000011",
      "100101111001" when "10110000100",
      "100101111000" when "10110000101",
      "100101111000" when "10110000110",
      "100101110111" when "10110000111",
      "100101110110" when "10110001000",
      "100101110101" when "10110001001",
      "100101110101" when "10110001010",
      "100101110100" when "10110001011",
      "100101110011" when "10110001100",
      "100101110011" when "10110001101",
      "100101110010" when "10110001110",
      "100101110001" when "10110001111",
      "100101110001" when "10110010000",
      "100101110000" when "10110010001",
      "100101101111" when "10110010010",
      "100101101110" when "10110010011",
      "100101101110" when "10110010100",
      "100101101101" when "10110010101",
      "100101101100" when "10110010110",
      "100101101100" when "10110010111",
      "100101101011" when "10110011000",
      "100101101010" when "10110011001",
      "100101101010" when "10110011010",
      "100101101001" when "10110011011",
      "100101101000" when "10110011100",
      "100101101000" when "10110011101",
      "100101100111" when "10110011110",
      "100101100110" when "10110011111",
      "100101100101" when "10110100000",
      "100101100101" when "10110100001",
      "100101100100" when "10110100010",
      "100101100011" when "10110100011",
      "100101100011" when "10110100100",
      "100101100010" when "10110100101",
      "100101100001" when "10110100110",
      "100101100001" when "10110100111",
      "100101100000" when "10110101000",
      "100101011111" when "10110101001",
      "100101011111" when "10110101010",
      "100101011110" when "10110101011",
      "100101011101" when "10110101100",
      "100101011101" when "10110101101",
      "100101011100" when "10110101110",
      "100101011011" when "10110101111",
      "100101011011" when "10110110000",
      "100101011010" when "10110110001",
      "100101011001" when "10110110010",
      "100101011000" when "10110110011",
      "100101011000" when "10110110100",
      "100101010111" when "10110110101",
      "100101010110" when "10110110110",
      "100101010110" when "10110110111",
      "100101010101" when "10110111000",
      "100101010100" when "10110111001",
      "100101010100" when "10110111010",
      "100101010011" when "10110111011",
      "100101010010" when "10110111100",
      "100101010010" when "10110111101",
      "100101010001" when "10110111110",
      "100101010000" when "10110111111",
      "100101010000" when "10111000000",
      "100101001111" when "10111000001",
      "100101001110" when "10111000010",
      "100101001110" when "10111000011",
      "100101001101" when "10111000100",
      "100101001100" when "10111000101",
      "100101001100" when "10111000110",
      "100101001011" when "10111000111",
      "100101001010" when "10111001000",
      "100101001010" when "10111001001",
      "100101001001" when "10111001010",
      "100101001000" when "10111001011",
      "100101001000" when "10111001100",
      "100101000111" when "10111001101",
      "100101000110" when "10111001110",
      "100101000110" when "10111001111",
      "100101000101" when "10111010000",
      "100101000100" when "10111010001",
      "100101000100" when "10111010010",
      "100101000011" when "10111010011",
      "100101000010" when "10111010100",
      "100101000001" when "10111010101",
      "100101000001" when "10111010110",
      "100101000000" when "10111010111",
      "100100111111" when "10111011000",
      "100100111111" when "10111011001",
      "100100111110" when "10111011010",
      "100100111101" when "10111011011",
      "100100111101" when "10111011100",
      "100100111100" when "10111011101",
      "100100111011" when "10111011110",
      "100100111011" when "10111011111",
      "100100111010" when "10111100000",
      "100100111001" when "10111100001",
      "100100111001" when "10111100010",
      "100100111000" when "10111100011",
      "100100111000" when "10111100100",
      "100100110111" when "10111100101",
      "100100110110" when "10111100110",
      "100100110110" when "10111100111",
      "100100110101" when "10111101000",
      "100100110100" when "10111101001",
      "100100110100" when "10111101010",
      "100100110011" when "10111101011",
      "100100110010" when "10111101100",
      "100100110010" when "10111101101",
      "100100110001" when "10111101110",
      "100100110000" when "10111101111",
      "100100110000" when "10111110000",
      "100100101111" when "10111110001",
      "100100101110" when "10111110010",
      "100100101110" when "10111110011",
      "100100101101" when "10111110100",
      "100100101100" when "10111110101",
      "100100101100" when "10111110110",
      "100100101011" when "10111110111",
      "100100101010" when "10111111000",
      "100100101010" when "10111111001",
      "100100101001" when "10111111010",
      "100100101000" when "10111111011",
      "100100101000" when "10111111100",
      "100100100111" when "10111111101",
      "100100100110" when "10111111110",
      "100100100110" when "10111111111",
      "100100100101" when "11000000000",
      "100100100100" when "11000000001",
      "100100100100" when "11000000010",
      "100100100011" when "11000000011",
      "100100100010" when "11000000100",
      "100100100010" when "11000000101",
      "100100100001" when "11000000110",
      "100100100001" when "11000000111",
      "100100100000" when "11000001000",
      "100100011111" when "11000001001",
      "100100011111" when "11000001010",
      "100100011110" when "11000001011",
      "100100011101" when "11000001100",
      "100100011101" when "11000001101",
      "100100011100" when "11000001110",
      "100100011011" when "11000001111",
      "100100011011" when "11000010000",
      "100100011010" when "11000010001",
      "100100011001" when "11000010010",
      "100100011001" when "11000010011",
      "100100011000" when "11000010100",
      "100100010111" when "11000010101",
      "100100010111" when "11000010110",
      "100100010110" when "11000010111",
      "100100010110" when "11000011000",
      "100100010101" when "11000011001",
      "100100010100" when "11000011010",
      "100100010100" when "11000011011",
      "100100010011" when "11000011100",
      "100100010010" when "11000011101",
      "100100010010" when "11000011110",
      "100100010001" when "11000011111",
      "100100010000" when "11000100000",
      "100100010000" when "11000100001",
      "100100001111" when "11000100010",
      "100100001110" when "11000100011",
      "100100001110" when "11000100100",
      "100100001101" when "11000100101",
      "100100001101" when "11000100110",
      "100100001100" when "11000100111",
      "100100001011" when "11000101000",
      "100100001011" when "11000101001",
      "100100001010" when "11000101010",
      "100100001001" when "11000101011",
      "100100001001" when "11000101100",
      "100100001000" when "11000101101",
      "100100000111" when "11000101110",
      "100100000111" when "11000101111",
      "100100000110" when "11000110000",
      "100100000110" when "11000110001",
      "100100000101" when "11000110010",
      "100100000100" when "11000110011",
      "100100000100" when "11000110100",
      "100100000011" when "11000110101",
      "100100000010" when "11000110110",
      "100100000010" when "11000110111",
      "100100000001" when "11000111000",
      "100100000000" when "11000111001",
      "100100000000" when "11000111010",
      "100011111111" when "11000111011",
      "100011111111" when "11000111100",
      "100011111110" when "11000111101",
      "100011111101" when "11000111110",
      "100011111101" when "11000111111",
      "100011111100" when "11001000000",
      "100011111011" when "11001000001",
      "100011111011" when "11001000010",
      "100011111010" when "11001000011",
      "100011111001" when "11001000100",
      "100011111001" when "11001000101",
      "100011111000" when "11001000110",
      "100011111000" when "11001000111",
      "100011110111" when "11001001000",
      "100011110110" when "11001001001",
      "100011110110" when "11001001010",
      "100011110101" when "11001001011",
      "100011110100" when "11001001100",
      "100011110100" when "11001001101",
      "100011110011" when "11001001110",
      "100011110011" when "11001001111",
      "100011110010" when "11001010000",
      "100011110001" when "11001010001",
      "100011110001" when "11001010010",
      "100011110000" when "11001010011",
      "100011101111" when "11001010100",
      "100011101111" when "11001010101",
      "100011101110" when "11001010110",
      "100011101110" when "11001010111",
      "100011101101" when "11001011000",
      "100011101100" when "11001011001",
      "100011101100" when "11001011010",
      "100011101011" when "11001011011",
      "100011101010" when "11001011100",
      "100011101010" when "11001011101",
      "100011101001" when "11001011110",
      "100011101001" when "11001011111",
      "100011101000" when "11001100000",
      "100011100111" when "11001100001",
      "100011100111" when "11001100010",
      "100011100110" when "11001100011",
      "100011100110" when "11001100100",
      "100011100101" when "11001100101",
      "100011100100" when "11001100110",
      "100011100100" when "11001100111",
      "100011100011" when "11001101000",
      "100011100010" when "11001101001",
      "100011100010" when "11001101010",
      "100011100001" when "11001101011",
      "100011100001" when "11001101100",
      "100011100000" when "11001101101",
      "100011011111" when "11001101110",
      "100011011111" when "11001101111",
      "100011011110" when "11001110000",
      "100011011110" when "11001110001",
      "100011011101" when "11001110010",
      "100011011100" when "11001110011",
      "100011011100" when "11001110100",
      "100011011011" when "11001110101",
      "100011011010" when "11001110110",
      "100011011010" when "11001110111",
      "100011011001" when "11001111000",
      "100011011001" when "11001111001",
      "100011011000" when "11001111010",
      "100011010111" when "11001111011",
      "100011010111" when "11001111100",
      "100011010110" when "11001111101",
      "100011010110" when "11001111110",
      "100011010101" when "11001111111",
      "100011010100" when "11010000000",
      "100011010100" when "11010000001",
      "100011010011" when "11010000010",
      "100011010011" when "11010000011",
      "100011010010" when "11010000100",
      "100011010001" when "11010000101",
      "100011010001" when "11010000110",
      "100011010000" when "11010000111",
      "100011010000" when "11010001000",
      "100011001111" when "11010001001",
      "100011001110" when "11010001010",
      "100011001110" when "11010001011",
      "100011001101" when "11010001100",
      "100011001100" when "11010001101",
      "100011001100" when "11010001110",
      "100011001011" when "11010001111",
      "100011001011" when "11010010000",
      "100011001010" when "11010010001",
      "100011001001" when "11010010010",
      "100011001001" when "11010010011",
      "100011001000" when "11010010100",
      "100011001000" when "11010010101",
      "100011000111" when "11010010110",
      "100011000110" when "11010010111",
      "100011000110" when "11010011000",
      "100011000101" when "11010011001",
      "100011000101" when "11010011010",
      "100011000100" when "11010011011",
      "100011000011" when "11010011100",
      "100011000011" when "11010011101",
      "100011000010" when "11010011110",
      "100011000010" when "11010011111",
      "100011000001" when "11010100000",
      "100011000000" when "11010100001",
      "100011000000" when "11010100010",
      "100010111111" when "11010100011",
      "100010111111" when "11010100100",
      "100010111110" when "11010100101",
      "100010111101" when "11010100110",
      "100010111101" when "11010100111",
      "100010111100" when "11010101000",
      "100010111100" when "11010101001",
      "100010111011" when "11010101010",
      "100010111010" when "11010101011",
      "100010111010" when "11010101100",
      "100010111001" when "11010101101",
      "100010111001" when "11010101110",
      "100010111000" when "11010101111",
      "100010111000" when "11010110000",
      "100010110111" when "11010110001",
      "100010110110" when "11010110010",
      "100010110110" when "11010110011",
      "100010110101" when "11010110100",
      "100010110101" when "11010110101",
      "100010110100" when "11010110110",
      "100010110011" when "11010110111",
      "100010110011" when "11010111000",
      "100010110010" when "11010111001",
      "100010110010" when "11010111010",
      "100010110001" when "11010111011",
      "100010110000" when "11010111100",
      "100010110000" when "11010111101",
      "100010101111" when "11010111110",
      "100010101111" when "11010111111",
      "100010101110" when "11011000000",
      "100010101101" when "11011000001",
      "100010101101" when "11011000010",
      "100010101100" when "11011000011",
      "100010101100" when "11011000100",
      "100010101011" when "11011000101",
      "100010101011" when "11011000110",
      "100010101010" when "11011000111",
      "100010101001" when "11011001000",
      "100010101001" when "11011001001",
      "100010101000" when "11011001010",
      "100010101000" when "11011001011",
      "100010100111" when "11011001100",
      "100010100110" when "11011001101",
      "100010100110" when "11011001110",
      "100010100101" when "11011001111",
      "100010100101" when "11011010000",
      "100010100100" when "11011010001",
      "100010100100" when "11011010010",
      "100010100011" when "11011010011",
      "100010100010" when "11011010100",
      "100010100010" when "11011010101",
      "100010100001" when "11011010110",
      "100010100001" when "11011010111",
      "100010100000" when "11011011000",
      "100010011111" when "11011011001",
      "100010011111" when "11011011010",
      "100010011110" when "11011011011",
      "100010011110" when "11011011100",
      "100010011101" when "11011011101",
      "100010011101" when "11011011110",
      "100010011100" when "11011011111",
      "100010011011" when "11011100000",
      "100010011011" when "11011100001",
      "100010011010" when "11011100010",
      "100010011010" when "11011100011",
      "100010011001" when "11011100100",
      "100010011001" when "11011100101",
      "100010011000" when "11011100110",
      "100010010111" when "11011100111",
      "100010010111" when "11011101000",
      "100010010110" when "11011101001",
      "100010010110" when "11011101010",
      "100010010101" when "11011101011",
      "100010010100" when "11011101100",
      "100010010100" when "11011101101",
      "100010010011" when "11011101110",
      "100010010011" when "11011101111",
      "100010010010" when "11011110000",
      "100010010010" when "11011110001",
      "100010010001" when "11011110010",
      "100010010000" when "11011110011",
      "100010010000" when "11011110100",
      "100010001111" when "11011110101",
      "100010001111" when "11011110110",
      "100010001110" when "11011110111",
      "100010001110" when "11011111000",
      "100010001101" when "11011111001",
      "100010001100" when "11011111010",
      "100010001100" when "11011111011",
      "100010001011" when "11011111100",
      "100010001011" when "11011111101",
      "100010001010" when "11011111110",
      "100010001010" when "11011111111",
      "100010001001" when "11100000000",
      "100010001000" when "11100000001",
      "100010001000" when "11100000010",
      "100010000111" when "11100000011",
      "100010000111" when "11100000100",
      "100010000110" when "11100000101",
      "100010000110" when "11100000110",
      "100010000101" when "11100000111",
      "100010000100" when "11100001000",
      "100010000100" when "11100001001",
      "100010000011" when "11100001010",
      "100010000011" when "11100001011",
      "100010000010" when "11100001100",
      "100010000010" when "11100001101",
      "100010000001" when "11100001110",
      "100010000001" when "11100001111",
      "100010000000" when "11100010000",
      "100001111111" when "11100010001",
      "100001111111" when "11100010010",
      "100001111110" when "11100010011",
      "100001111110" when "11100010100",
      "100001111101" when "11100010101",
      "100001111101" when "11100010110",
      "100001111100" when "11100010111",
      "100001111011" when "11100011000",
      "100001111011" when "11100011001",
      "100001111010" when "11100011010",
      "100001111010" when "11100011011",
      "100001111001" when "11100011100",
      "100001111001" when "11100011101",
      "100001111000" when "11100011110",
      "100001111000" when "11100011111",
      "100001110111" when "11100100000",
      "100001110110" when "11100100001",
      "100001110110" when "11100100010",
      "100001110101" when "11100100011",
      "100001110101" when "11100100100",
      "100001110100" when "11100100101",
      "100001110100" when "11100100110",
      "100001110011" when "11100100111",
      "100001110011" when "11100101000",
      "100001110010" when "11100101001",
      "100001110001" when "11100101010",
      "100001110001" when "11100101011",
      "100001110000" when "11100101100",
      "100001110000" when "11100101101",
      "100001101111" when "11100101110",
      "100001101111" when "11100101111",
      "100001101110" when "11100110000",
      "100001101110" when "11100110001",
      "100001101101" when "11100110010",
      "100001101100" when "11100110011",
      "100001101100" when "11100110100",
      "100001101011" when "11100110101",
      "100001101011" when "11100110110",
      "100001101010" when "11100110111",
      "100001101010" when "11100111000",
      "100001101001" when "11100111001",
      "100001101001" when "11100111010",
      "100001101000" when "11100111011",
      "100001100111" when "11100111100",
      "100001100111" when "11100111101",
      "100001100110" when "11100111110",
      "100001100110" when "11100111111",
      "100001100101" when "11101000000",
      "100001100101" when "11101000001",
      "100001100100" when "11101000010",
      "100001100100" when "11101000011",
      "100001100011" when "11101000100",
      "100001100010" when "11101000101",
      "100001100010" when "11101000110",
      "100001100001" when "11101000111",
      "100001100001" when "11101001000",
      "100001100000" when "11101001001",
      "100001100000" when "11101001010",
      "100001011111" when "11101001011",
      "100001011111" when "11101001100",
      "100001011110" when "11101001101",
      "100001011110" when "11101001110",
      "100001011101" when "11101001111",
      "100001011100" when "11101010000",
      "100001011100" when "11101010001",
      "100001011011" when "11101010010",
      "100001011011" when "11101010011",
      "100001011010" when "11101010100",
      "100001011010" when "11101010101",
      "100001011001" when "11101010110",
      "100001011001" when "11101010111",
      "100001011000" when "11101011000",
      "100001011000" when "11101011001",
      "100001010111" when "11101011010",
      "100001010110" when "11101011011",
      "100001010110" when "11101011100",
      "100001010101" when "11101011101",
      "100001010101" when "11101011110",
      "100001010100" when "11101011111",
      "100001010100" when "11101100000",
      "100001010011" when "11101100001",
      "100001010011" when "11101100010",
      "100001010010" when "11101100011",
      "100001010010" when "11101100100",
      "100001010001" when "11101100101",
      "100001010001" when "11101100110",
      "100001010000" when "11101100111",
      "100001001111" when "11101101000",
      "100001001111" when "11101101001",
      "100001001110" when "11101101010",
      "100001001110" when "11101101011",
      "100001001101" when "11101101100",
      "100001001101" when "11101101101",
      "100001001100" when "11101101110",
      "100001001100" when "11101101111",
      "100001001011" when "11101110000",
      "100001001011" when "11101110001",
      "100001001010" when "11101110010",
      "100001001010" when "11101110011",
      "100001001001" when "11101110100",
      "100001001000" when "11101110101",
      "100001001000" when "11101110110",
      "100001000111" when "11101110111",
      "100001000111" when "11101111000",
      "100001000110" when "11101111001",
      "100001000110" when "11101111010",
      "100001000101" when "11101111011",
      "100001000101" when "11101111100",
      "100001000100" when "11101111101",
      "100001000100" when "11101111110",
      "100001000011" when "11101111111",
      "100001000011" when "11110000000",
      "100001000010" when "11110000001",
      "100001000001" when "11110000010",
      "100001000001" when "11110000011",
      "100001000000" when "11110000100",
      "100001000000" when "11110000101",
      "100000111111" when "11110000110",
      "100000111111" when "11110000111",
      "100000111110" when "11110001000",
      "100000111110" when "11110001001",
      "100000111101" when "11110001010",
      "100000111101" when "11110001011",
      "100000111100" when "11110001100",
      "100000111100" when "11110001101",
      "100000111011" when "11110001110",
      "100000111011" when "11110001111",
      "100000111010" when "11110010000",
      "100000111010" when "11110010001",
      "100000111001" when "11110010010",
      "100000111000" when "11110010011",
      "100000111000" when "11110010100",
      "100000110111" when "11110010101",
      "100000110111" when "11110010110",
      "100000110110" when "11110010111",
      "100000110110" when "11110011000",
      "100000110101" when "11110011001",
      "100000110101" when "11110011010",
      "100000110100" when "11110011011",
      "100000110100" when "11110011100",
      "100000110011" when "11110011101",
      "100000110011" when "11110011110",
      "100000110010" when "11110011111",
      "100000110010" when "11110100000",
      "100000110001" when "11110100001",
      "100000110001" when "11110100010",
      "100000110000" when "11110100011",
      "100000110000" when "11110100100",
      "100000101111" when "11110100101",
      "100000101111" when "11110100110",
      "100000101110" when "11110100111",
      "100000101101" when "11110101000",
      "100000101101" when "11110101001",
      "100000101100" when "11110101010",
      "100000101100" when "11110101011",
      "100000101011" when "11110101100",
      "100000101011" when "11110101101",
      "100000101010" when "11110101110",
      "100000101010" when "11110101111",
      "100000101001" when "11110110000",
      "100000101001" when "11110110001",
      "100000101000" when "11110110010",
      "100000101000" when "11110110011",
      "100000100111" when "11110110100",
      "100000100111" when "11110110101",
      "100000100110" when "11110110110",
      "100000100110" when "11110110111",
      "100000100101" when "11110111000",
      "100000100101" when "11110111001",
      "100000100100" when "11110111010",
      "100000100100" when "11110111011",
      "100000100011" when "11110111100",
      "100000100011" when "11110111101",
      "100000100010" when "11110111110",
      "100000100010" when "11110111111",
      "100000100001" when "11111000000",
      "100000100000" when "11111000001",
      "100000100000" when "11111000010",
      "100000011111" when "11111000011",
      "100000011111" when "11111000100",
      "100000011110" when "11111000101",
      "100000011110" when "11111000110",
      "100000011101" when "11111000111",
      "100000011101" when "11111001000",
      "100000011100" when "11111001001",
      "100000011100" when "11111001010",
      "100000011011" when "11111001011",
      "100000011011" when "11111001100",
      "100000011010" when "11111001101",
      "100000011010" when "11111001110",
      "100000011001" when "11111001111",
      "100000011001" when "11111010000",
      "100000011000" when "11111010001",
      "100000011000" when "11111010010",
      "100000010111" when "11111010011",
      "100000010111" when "11111010100",
      "100000010110" when "11111010101",
      "100000010110" when "11111010110",
      "100000010101" when "11111010111",
      "100000010101" when "11111011000",
      "100000010100" when "11111011001",
      "100000010100" when "11111011010",
      "100000010011" when "11111011011",
      "100000010011" when "11111011100",
      "100000010010" when "11111011101",
      "100000010010" when "11111011110",
      "100000010001" when "11111011111",
      "100000010001" when "11111100000",
      "100000010000" when "11111100001",
      "100000010000" when "11111100010",
      "100000001111" when "11111100011",
      "100000001111" when "11111100100",
      "100000001110" when "11111100101",
      "100000001110" when "11111100110",
      "100000001101" when "11111100111",
      "100000001101" when "11111101000",
      "100000001100" when "11111101001",
      "100000001100" when "11111101010",
      "100000001011" when "11111101011",
      "100000001011" when "11111101100",
      "100000001010" when "11111101101",
      "100000001010" when "11111101110",
      "100000001001" when "11111101111",
      "100000001001" when "11111110000",
      "100000001000" when "11111110001",
      "100000001000" when "11111110010",
      "100000000111" when "11111110011",
      "100000000111" when "11111110100",
      "100000000110" when "11111110101",
      "100000000110" when "11111110110",
      "100000000101" when "11111110111",
      "100000000101" when "11111111000",
      "100000000100" when "11111111001",
      "100000000100" when "11111111010",
      "100000000011" when "11111111011",
      "100000000011" when "11111111100",
      "100000000010" when "11111111101",
      "100000000010" when "11111111110",
      "100000000001" when "11111111111",
      "------------" when others;
   Y1_c0 <= Y0_c0; -- for the possible blockram register
   Y <= Y1_c0;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_80_Freq300_uid18
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_80_Freq300_uid18 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(79 downto 0);
          Y : in  std_logic_vector(79 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(79 downto 0)   );
end entity;

architecture arch of IntAdder_80_Freq300_uid18 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2 :  std_logic;
signal X_0_c1, X_0_c2 :  std_logic_vector(15 downto 0);
signal Y_0_c1, Y_0_c2 :  std_logic_vector(15 downto 0);
signal S_0_c2 :  std_logic_vector(15 downto 0);
signal R_0_c2 :  std_logic_vector(14 downto 0);
signal Cin_1_c2 :  std_logic;
signal X_1_c1, X_1_c2 :  std_logic_vector(65 downto 0);
signal Y_1_c1, Y_1_c2 :  std_logic_vector(65 downto 0);
signal S_1_c2 :  std_logic_vector(65 downto 0);
signal R_1_c2 :  std_logic_vector(64 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
               X_0_c2 <= X_0_c1;
               Y_0_c2 <= Y_0_c1;
               X_1_c2 <= X_1_c1;
               Y_1_c2 <= Y_1_c1;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c1 <= '0' & X(14 downto 0);
   Y_0_c1 <= '0' & Y(14 downto 0);
   S_0_c2 <= X_0_c2 + Y_0_c2 + Cin_0_c2;
   R_0_c2 <= S_0_c2(14 downto 0);
   Cin_1_c2 <= S_0_c2(15);
   X_1_c1 <= '0' & X(79 downto 15);
   Y_1_c1 <= '0' & Y(79 downto 15);
   S_1_c2 <= X_1_c2 + Y_1_c2 + Cin_1_c2;
   R_1_c2 <= S_1_c2(64 downto 0);
   R <= R_1_c2 & R_0_c2 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_80_Freq300_uid21
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_80_Freq300_uid21 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(79 downto 0);
          Y : in  std_logic_vector(79 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(79 downto 0)   );
end entity;

architecture arch of IntAdder_80_Freq300_uid21 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3 :  std_logic;
signal X_0_c2, X_0_c3 :  std_logic_vector(67 downto 0);
signal Y_0_c2, Y_0_c3 :  std_logic_vector(67 downto 0);
signal S_0_c3 :  std_logic_vector(67 downto 0);
signal R_0_c3 :  std_logic_vector(66 downto 0);
signal Cin_1_c3 :  std_logic;
signal X_1_c2, X_1_c3 :  std_logic_vector(13 downto 0);
signal Y_1_c2, Y_1_c3 :  std_logic_vector(13 downto 0);
signal S_1_c3 :  std_logic_vector(13 downto 0);
signal R_1_c3 :  std_logic_vector(12 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
               X_0_c3 <= X_0_c2;
               Y_0_c3 <= Y_0_c2;
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c2 <= '0' & X(66 downto 0);
   Y_0_c2 <= '0' & Y(66 downto 0);
   S_0_c3 <= X_0_c3 + Y_0_c3 + Cin_0_c3;
   R_0_c3 <= S_0_c3(66 downto 0);
   Cin_1_c3 <= S_0_c3(67);
   X_1_c2 <= '0' & X(79 downto 67);
   Y_1_c2 <= '0' & Y(79 downto 67);
   S_1_c3 <= X_1_c3 + Y_1_c3 + Cin_1_c3;
   R_1_c3 <= S_1_c3(12 downto 0);
   R <= R_1_c3 & R_0_c3 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_79_Freq300_uid24
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_79_Freq300_uid24 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(78 downto 0);
          Y : in  std_logic_vector(78 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(78 downto 0)   );
end entity;

architecture arch of IntAdder_79_Freq300_uid24 is
signal Rtmp_c4 :  std_logic_vector(78 downto 0);
signal X_c4 :  std_logic_vector(78 downto 0);
signal Y_c4 :  std_logic_vector(78 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               X_c4 <= X;
               Y_c4 <= Y;
               Cin_c4 <= Cin_c3;
            end if;
         end if;
      end process;
   Rtmp_c4 <= X_c4 + Y_c4 + Cin_c4;
   R <= Rtmp_c4;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_79_Freq300_uid27
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_79_Freq300_uid27 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(78 downto 0);
          Y : in  std_logic_vector(78 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(78 downto 0)   );
end entity;

architecture arch of IntAdder_79_Freq300_uid27 is
signal Rtmp_c5 :  std_logic_vector(78 downto 0);
signal X_c5 :  std_logic_vector(78 downto 0);
signal Y_c5 :  std_logic_vector(78 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               X_c5 <= X;
               Y_c5 <= Y;
               Cin_c5 <= Cin_c4;
            end if;
         end if;
      end process;
   Rtmp_c5 <= X_c5 + Y_c5 + Cin_c5;
   R <= Rtmp_c5;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_70_Freq300_uid30
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_70_Freq300_uid30 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(69 downto 0);
          Y : in  std_logic_vector(69 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(69 downto 0)   );
end entity;

architecture arch of IntAdder_70_Freq300_uid30 is
signal Rtmp_c5 :  std_logic_vector(69 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
         end if;
      end process;
   Rtmp_c5 <= X + Y + Cin_c5;
   R <= Rtmp_c5;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_70_Freq300_uid33
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_70_Freq300_uid33 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(69 downto 0);
          Y : in  std_logic_vector(69 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(69 downto 0)   );
end entity;

architecture arch of IntAdder_70_Freq300_uid33 is
signal Rtmp_c6 :  std_logic_vector(69 downto 0);
signal X_c6 :  std_logic_vector(69 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X;
               Cin_c6 <= Cin_c5;
            end if;
         end if;
      end process;
   Rtmp_c6 <= X_c6 + Y + Cin_c6;
   R <= Rtmp_c6;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_70_Freq300_uid36
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_70_Freq300_uid36 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7 : in std_logic;
          X : in  std_logic_vector(69 downto 0);
          Y : in  std_logic_vector(69 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(69 downto 0)   );
end entity;

architecture arch of IntAdder_70_Freq300_uid36 is
signal Rtmp_c7 :  std_logic_vector(69 downto 0);
signal X_c7 :  std_logic_vector(69 downto 0);
signal Y_c7 :  std_logic_vector(69 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               X_c7 <= X;
               Y_c7 <= Y;
               Cin_c7 <= Cin_c6;
            end if;
         end if;
      end process;
   Rtmp_c7 <= X_c7 + Y_c7 + Cin_c7;
   R <= Rtmp_c7;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable0_Freq300_uid38
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable0_Freq300_uid38 is
    port (clk : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : out  std_logic_vector(103 downto 0)   );
end entity;

architecture arch of LogTable0_Freq300_uid38 is
signal Y0_c0 :  std_logic_vector(103 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c0 :  std_logic_vector(103 downto 0);
begin
   with X  select  Y0_c0 <= 
      "11111111111111111011111111111111101111111111111111000000000000000000000000000000000000000000000000000000" when "00000000000",
      "11111111111111111011111111111111101111111111111111000000000000000000000000000000000000000000000000000000" when "00000000001",
      "00000000000111111100000111111111111010101010111001101011000100010001101110111100111000000110111000001000" when "00000000010",
      "00000000001111111100100000000001000101011001010100100010001001001100110101011111001101011111100001111101" when "00000000011",
      "00000000010111111101001000000100010000010100010000100001010100011001110011111001110101100001101111001011" when "00000000100",
      "00000000011111111110000000001010011011101010110000000100111011110011100000110011100011110111011101100000" when "00000000101",
      "00000000100111111111001000010100100111110001110111111001111000011011110110000100110111010010110111100111" when "00000000110",
      "00000000110000000000100000100011110101000100101111101110000000110100101101010011100001100000011000101000" when "00000000111",
      "00000000111000000010001000111001000100000100100011000000101010111110100110110001100011100101011001011101" when "00000001000",
      "00000001000000000100000001010101010101011000100001110011010101111110010110011000111000110011110110001110" when "00000001001",
      "00000001001000000110001001111001101001101110000001011010011011001011010010010001001110010011110101001110" when "00000001010",
      "00000001010000001000100010100111000001111000011101001110000111000111011111000001110000000000000001100010" when "00000001011",
      "00000001011000001011001011011110011110110001010111011011011010000011010110000100100010010001011101010011" when "00000001100",
      "00000001100000001110000100100001000001011000011001110101010000001110000010100101110011111100100110111100" when "00000001101",
      "00000001101000010001001101101111101010110011010110100101110001110100010010001101101101001110000100100101" when "00000001110",
      "00000001110000010100100111001011011100001110001000111111101010101110110110100111011110101001111110110011" when "00000001111",
      "00000001111000011000010000110101010110111010110110001111101010000010010101101101110110110000000100001010" when "00000010000",
      "00000010000000011100001010101110011100010001101110001110001001010001100110011000101101010000010111110100" when "00000010001",
      "00000010001000100000010100110111101101110001001100010000111011100100010111111101000001010011101100010000" when "00000010010",
      "00000010010000100100101111010010001100111101110111111101000100100011100011000100111010011111111110110011" when "00000010011",
      "00000010011000101001011001111110111011100010100101111000110111001100100010111010010101010110001111001110" when "00000010100",
      "00000010100000101110010100111110111011010000011000011101111100011101010101110100000001001101101000011111" when "00000010101",
      "00000010101000110011100000010011001101111110100000101011100001111010100101001001011000101000111100011010" when "00000010110",
      "00000010110000111000111011111100110101101010011110111000110000010001010100000111000101010000110010110100" when "00000010111",
      "00000010111000111110100111111100110100011000000011100111001001110101110101110011001110000000100000001000" when "00000011000",
      "00000011000001000100100100010100001100010001010000010101010001000001001011000101100001001101111111000010" when "00000011001",
      "00000011001001001010110001000011111111100110011000010001010110101110101001001101000100101000100111111011" when "00000011010",
      "00000011010001010001001110001101010000101110000001001100010000111011001010010010110010111000110111101110" when "00000011011",
      "00000011011001010111111011110001000010000101000100001100011001000111101001011101010001010100001011110011" when "00000011100",
      "00000011100001011110111001110000010110001110101110100000110011000000001100010000010001100000001001100001" when "00000011101",
      "00000011101001100110001000001100001111110100100010010100011011001001011011111000000000000101111101011001" when "00000011110",
      "00000011110001101101100111000101110001100110010111100001011101110101110000100101110101111110011000001111" when "00000011111",
      "00000011111001110101010110011101111110011010011100100100110110000011110010011010011010000111010111011000" when "00000100000",
      "00000100000001111101010110010101111001001101010111010001110100100111110010001110100001000001011011100111" when "00000100001",
      "00000100001010000101100110101110100101000010000101100101101111100001011111000010111011000100111111111101" when "00000100010",
      "00000100010010001110000111101001000101000001111110011011111001011111111011010100101100111001001010000010" when "00000100011",
      "00000100011010010110111001000110011100011100110010100001100001110100110110101010011100010110111010110011" when "00000100100",
      "00000100100010011111111011000111101110101000101101001001111100011001010000100100110010001111111100011111" when "00000100101",
      "00000100101010101001001101101101111111000010010101000010110010000100101001010011001011000111010011000101" when "00000100110",
      "00000100110010110010110000111010010001001100101101001000011001011000100110000100010010101111110111011110" when "00000100111",
      "00000100111010111100100100101101101000110001010101011010010111100010001110100000001011111000001010100010" when "00000101000",
      "00000101000011000110101001001001001001100000001011110000001001110011001001010000110001101111111110111110" when "00000101001",
      "00000101001011010000111110001101110111001111101100101101110111010011011110010100010011001011100000100010" when "00000101010",
      "00000101010011011011100011111100110101111100110100011001001011001110100101101011111110010010100110010110" when "00000101011",
      "00000101011011100110011010010111001001101010111111001110010111011100001001110000010001101011110001010110" when "00000101100",
      "00000101100011110001100001011101110110100100001010110101011111100111000100101011001011001010100000110110" when "00000101101",
      "00000101100011110001100001011101110110100100001010110101011111100111000100101011001011001010100000110110" when "00000101110",
      "00000101101011111100111001010010000000111000110110110111101100110100000000101111110101011001110010100011" when "00000101111",
      "00000101110100001000100001110100101101000000000101110100101001101001000011111110100101000111011110000100" when "00000110000",
      "00000101111100010100011011000110111111010111011101111000000110111000001111011011001011011101110010000000" when "00000110001",
      "00000110000100100000100101001001111100100011001001101111101000101110011011010010111110011110011000000110" when "00000110010",
      "00000110001100101100111111111110101001001101111001100000011100101000011001000111111001011000111100110111" when "00000110011",
      "00000110010100111001101011100110001010001001000011011101010111101111100101101100111101111111010100010110" when "00000110100",
      "00000110011101000110101000000001100100001100100100111100111110000000010100111000101101000100000111100001" when "00000110101",
      "00000110100101010011110101010001111100010111000011001111110001111011000001101001011111100001101101010000" when "00000110110",
      "00000110101101100001010011011000010111101101101100010110101101000010001101010000000010111101111110100111" when "00000110111",
      "00000110110101101111000010010101111011011100010111111001100001000110111000101011111011111111101000000110" when "00000111000",
      "00000110111101111101000010001011101100110101100111111101100010000101000011111110010110010011100101000100" when "00000111001",
      "00000111000110001011010010111010110001010010101001111100011000110001111111001111010110010111100101000010" when "00000111010",
      "00000111001110011001110100100100001110010011010111011010111110011101111001111010010010100011001100001011" when "00000111011",
      "00000111010110101000100111001001001001011110010111000000100001001010111100101110010001111100011110011011" when "00000111100",
      "00000111011110110111101010101010101000100000111101001101110000111010111011101000001101101011001000011100" when "00000111101",
      "00000111100111000110111111001001110001001111001101010100010101110101101101000100010110010101110010101011" when "00000111110",
      "00000111101111010110100100100111101001100011111010001110001111001001110100011110001010100011010001100111" when "00000111111",
      "00000111110111100110011011000101010111100000100111010101011011001001001110001101111100111110101110001001" when "00001000000",
      "00000111111111110110100010100100000001001101101001011011101000000011101011101100100000011011100000110101" when "00001000001",
      "00000111111111110110100010100100000001001101101001011011101000000011101011101100100000011011100000110101" when "00001000010",
      "00001000001000000110111011000100101100111010000111100010001110000000101110011110001110101110101001101100" when "00001000011",
      "00001000010000010111100100101000100000111011111011110010010001111010110010000000000100001000100001110100" when "00001000100",
      "00001000011000101000011111010000100011101111110100010100110001011101010011101001110100001101110110100010" when "00001000101",
      "00001000100000111001101010111101111011111001010100001010111000000111101001010010101111000010100110000011" when "00001000110",
      "00001000101001001011000111110001110000000010110100000110011101010110010110111110100101110000001100010100" when "00001000111",
      "00001000110001011100110101101101000110111101100011100010101011110100110100110010111100101010101111111111" when "00001001000",
      "00001000111001101110110100110001000111100001101001011100110001111000110110001101111110011001100010010100" when "00001001001",
      "00001001000010000001000100111110111000101110000101001100111011001010000100110001101111101111100111000111" when "00001001010",
      "00001001001010010011100110010111100001101000101111011111010011010111000000010000110110110011110101001110" when "00001001011",
      "00001001010010100110011000111100001001011110011011001101010010011001010111000011000001010101110001101011" when "00001001100",
      "00001001011010111001011100101101110111100010110110010110110001101011101001100010010110011001001011111000" when "00001001101",
      "00001001100011001100110001101101110011010000101010111011101010110001101100001100000110011101010101101110" when "00001001110",
      "00001001101011100000010111111101000100001001011111110101011111010101111011111001111010110011010101011000" when "00001001111",
      "00001001101011100000010111111101000100001001011111110101011111010101111011111001111010110011010101011000" when "00001010000",
      "00001001110011110100001111011100110001110101111001110001001010011101011001000010111001010111011101111111" when "00001010001",
      "00001001111100001000011000001110000100000101011100001000111011010011111101101110001101111000111001001000" when "00001010010",
      "00001010000100011100110010010010000010101110101001111110011001010011000100011011101011001001010010110001" when "00001010011",
      "00001010001100110001011101101001110101101111000110110100110001100100010100100001000000010110101111011001" when "00001010100",
      "00001010010101000110011010010110100101001011010111101011001110000010001010010101101110110101110111101010" when "00001010101",
      "00001010011101011011101000011001011001001111000011110111010101111000010001100010000011000100011001001010" when "00001010110",
      "00001010100101110001000111110011011010001100110101111111110111100101101000000000010010001101100010101000" when "00001010111",
      "00001010101110000110111000100101110000011110011100110111011100100010000000111011100010011101011111110010" when "00001011000",
      "00001010110110011100111010110001100100100100101100010111100110001000111111010001010000011000001111111010" when "00001011001",
      "00001010111110110011001110010111111111000111011110011011110100101011111111110110110110110101101000111101" when "00001011010",
      "00001011000111001001110011011010001000110101110011111100110111101101101011011111111001011001110011010110" when "00001011011",
      "00001011001111100000101001111001001010100101110101101100001000001000001001111100110010100000101111001100" when "00001011100",
      "00001011001111100000101001111001001010100101110101101100001000001000001001111100110010100000101111001100" when "00001011101",
      "00001011010111110111110001110110001101010100110101001111001100000000001111000101101111011111101000111110" when "00001011110",
      "00001011100000001111001011010010011010000111001101111011100100000111011100000001010100011000110001100110" when "00001011111",
      "00001011101000100110110110001110111010001000100101110010100011001110101110010001111000101001011011010101" when "00001100000",
      "00001011110000111110110010101100110110101011101110011101001111001011110111110001001100010110110011110010" when "00001100001",
      "00001011111001010111000000101101011001001010100110001000101011110011011010011101011011010000111100111111" when "00001100010",
      "00001100000001101111100000010001101011000110011000100010001111101001000011010111010000001011101100011100" when "00001100011",
      "00001100001010001000010001011010110110000111011111110100000010101000100000101100101111110000000101010011" when "00001100100",
      "00001100010010100001010100001010000011111101100101100001100110101000101111101001011101100110000010100010" when "00001100101",
      "00001100011010111010101000100000011110011111100011100100101001111011011110100000100010010001000101100110" when "00001100110",
      "00001100100011010100001110011111001111101011100101001010000011101011000000100010010011010101101010010100" when "00001100111",
      "00001100100011010100001110011111001111101011100101001010000011101011000000100010010011010101101010010100" when "00001101000",
      "00001100101011101110000110000111100001100111000111101110111010011000010001001011110001011001000110100010" when "00001101001",
      "00001100110100001000001111011010011110011110111011111101110100011011000100111011001001101111001010011001" when "00001101010",
      "00001100111100100010101010011001010000100111000110101100010010100110100110010001101011001110111100011100" when "00001101011",
      "00001101000100111101010111000101000010011011000001111000010100110011111110001000000110111000111010110110" when "00001101100",
      "00001101001101011000010101011110111110011101011101100110001000110101000110111000100101110010010000010110" when "00001101101",
      "00001101010101110011100101101000001111011000100000111110000011010001101010011101110110100001011100000101" when "00001101110",
      "00001101011110001111000111100001111111111101101011001010100010110000001011100101010100101111010110101000" when "00001101111",
      "00001101100110101010111011001101011011000101110100010110011101001101011011001111010101011000111001000011" when "00001110000",
      "00001101101111000111000000101011101011110001001110101011010111100011111011110110010010011010000111101011" when "00001110001",
      "00001101101111000111000000101011101011110001001110101011010111100011111011110110010010011010000111101011" when "00001110010",
      "00001101110111100011010111111101111101000111100111010000000111100101110011110011101000001111010101101111" when "00001110011",
      "00001110000000000000000001000101011010011000000111000111100000001010110001110111010111010100010110111000" when "00001110100",
      "00001110001000011100111100000011001110111001010100001111000111110100100110000101000011010001010101001011" when "00001110101",
      "00001110010000111010001000111000100110001001010010011110011001101011110010100111011001001000111100101110" when "00001110110",
      "00001110011001010111100111100110101011101101100100100101110000110110111000001001111101011111111000100000" when "00001110111",
      "00001110100001110101011000001110101011010011001101001101111110001110000010000111000010111011101111100101" when "00001111000",
      "00001110101010010011011010110001110000101110101111110111101000101101010111010110010001000010100110010010" when "00001111001",
      "00001110110010110001101111010001000111111100010001111010111000000111110100100111010011110101110111101101" when "00001111010",
      "00001110111011010000010101101101111100111111011011100111001010011100110110010011000011011110100010011001" when "00001111011",
      "00001110111011010000010101101101111100111111011011100111001010011100110110010011000011011110100010011001" when "00001111100",
      "00001111000011101111001110001001011100000011011001000011010011110010110111101100010100000111011010110000" when "00001111101",
      "00001111001100001110011000100100110001011010111011001101101000111000101110011000100110010111011100110001" when "00001111110",
      "00001111010100101101110101000001001001100000011000111100010100010000001000111000100001000011100110110101" when "00001111111",
      "00001111011101001101100011011111110000110101101111111101110110000011011000000110110110001001000010010011" when "00010000000",
      "00001111100101101101100100000001110100000100100101111001101110101000001011110100110101101110011111101010" when "00010000001",
      "00001111101110001101110110101000011111111110001001010001010011110010001010101001111011110010110101001110" when "00010000010",
      "00001111110110101110011011010101000001011011010010100000110000110110101110101100110111001111011111111001" when "00010000011",
      "00001111111111001111010010001000100101011100100101000000010001100100110000011100000011010100011110100010" when "00010000100",
      "00001111111111001111010010001000100101011100100101000000010001100100110000011100000011010100011110100010" when "00010000101",
      "00010000000111110000011011000100011001001010010000000101010111110010001001111011001111100001000100101110" when "00010000110",
      "00010000010000010001110110001001101001110100010000000100011100000001011100111100011101011101010011011000" when "00010000111",
      "00010000011000110011100011011001100100110010001111010010011001000001100111001010110000011100101000111100" when "00010001000",
      "00010000100001010101100010110101010111100011100111000110100010001010001111111101100110111111010100000011" when "00010001001",
      "00010000101001110111110100011110001111101111100000111100100100110110011011111100011011111101101000011110" when "00010001010",
      "00010000110010011010011000010101011011000100110111010110110101000000010010111010011011001011101100010011" when "00010001011",
      "00010000111010111101001110011100000111011010010111000000100100011111100101010011101011110101110011001001" when "00010001100",
      "00010000111010111101001110011100000111011010010111000000100100011111100101010011101011110101110011001001" when "00010001101",
      "00010001000011100000010110110011100010101110011111110000100101101101011110110101110010111001101101100110" when "00010001110",
      "00010001001100000011110001011100111011000111100101101011111001001111110100011110110111111000111101000110" when "00010001111",
      "00010001010100100111011110011001011110110011110010001000100110101101111100011111100111101111101011011110" when "00010010000",
      "00010001011101001011011101101010011100001001000100110001000000110001011111101110001011100100100000111000" when "00010010001",
      "00010001100101101111101111010001000001100101010100100110110100010101010011111001001100001011001010100110" when "00010010010",
      "00010001101110010100010011001110011101101110010001000110100011000100101111001100000111011000000001011010" when "00010010011",
      "00010001110110111001001001100011111111010001100011001011001001001101100101110111110001001001001111111000" when "00010010100",
      "00010001110110111001001001100011111111010001100011001011001001001101100101110111110001001001001111111000" when "00010010101",
      "00010001111111011110010010010010110101000100101110010001101110100111000011010011111000110100101011110100" when "00010010110",
      "00010010001000000011101101011100001110000101010001011101100011001111110000010000110001111011111011000101" when "00010010111",
      "00010010010000101001011011000001011001011000101000011100000111000101011000110010010000100100000001110111" when "00010011000",
      "00010010011001001111011011000011100110001100001100101001011101011000000100101111100010110111010001011100" when "00010011001",
      "00010010100001110101101101100100000011110101010110010100101011011011110110010110010100001111101011110111" when "00010011010",
      "00010010101010011100010010100100000001110001011101100100100010111010100010110001110010110100000101110000" when "00010011011",
      "00010010101010011100010010100100000001110001011101100100100010111010100010110001110010110100000101110000" when "00010011100",
      "00010010110011000011001010000100101111100101111011011100010111101000011001011001100101010001001111100010" when "00010011101",
      "00010010111011101010010100000111011101000000001011000001000000111101101110101110111110010000101111110110" when "00010011110",
      "00010011000100010001110000101101011001110101101010011110000110111000000000110010100010100010001111001000" when "00010011111",
      "00010011001100111001011111110111110110000011111100001011011010100100101010111111001000111011110111000011" when "00010100000",
      "00010011010101100001100001101000000001110000100111110010011010111000000000011010110110101000001111101010" when "00010100001",
      "00010011011110001001110101111111001101001001011011010100000100010010100011110001111110101100101000001011" when "00010100010",
      "00010011011110001001110101111111001101001001011011010100000100010010100011110001111110101100101000001011" when "00010100011",
      "00010011100110110010011100111110101000100100001100001110101100110111010100110011111010101100110011100111" when "00010100100",
      "00010011101111011011010110100111100100011110111000100100001011110101001011101101101001110110101101101001" when "00010100101",
      "00010011111000000100100010111011010001011111101000000000001101000101111011100001100110001111110011100110" when "00010100110",
      "00010100000000101110000001111011000000010100101100111110110000100101010101000000101010111101111111111010" when "00010100111",
      "00010100001001010111110011101000000001110100100101110010110101100010100100001100111011010111011110001010" when "00010101000",
      "00010100010010000001111000000011100110111101111101101101010001101110100011010010011010101011011011110010" when "00010101001",
      "00010100010010000001111000000011100110111101111101101101010001101110100011010010011010101011011011110010" when "00010101010",
      "00010100011010101100001111001111000000110111101110000011110100101001011110000111101100010100101100001110" when "00010101011",
      "00010100100011010110111001001011100000110000111111011000010110110010000010001100001000000000101111101010" when "00010101100",
      "00010100101100000001110101111010011000000001001010100000010100111000110111011111001001101110001010010101" when "00010101101",
      "00010100110100101101000101011100111000000111111001101100010111011010011111010000101100011110000100001011" when "00010101110",
      "00010100111101011000100111110100010010101101001001110000000110000010010110010000001111110001111110011111" when "00010101111",
      "00010101000110000100011101000001111001100001001011001010000111011001011000100101100010110011110110001010" when "00010110000",
      "00010101000110000100011101000001111001100001001011001010000111011001011000100101100010110011110110001010" when "00010110001",
      "00010101001110110000100101000110111110011100100011001100001101000010100110000011010101010101001001011110" when "00010110010",
      "00010101010111011101000000000100110011100000001101000011101011101000000110001010011110001110010111010000" when "00010110011",
      "00010101100000001001101101111100101010110101011011000001111111011011001011111001100000110101010011001110" when "00010110100",
      "00010101101000110110101110101111110110101101110111100101011101001001111001101010111110100001011111101011" when "00010110101",
      "00010101110001100100000010011111101001100011100110100010001111001100100110101010110000001101101011010001" when "00010110110",
      "00010101110001100100000010011111101001100011100110100010001111001100100110101010110000001101101011010001" when "00010110111",
      "00010101111010010001101001001101010101111001000110001011011111001110000111010001011100010111000100010100" when "00010111000",
      "00010110000010111111100010111010001110011001010000011100101100010000111010111011000001001010010101111001" when "00010111001",
      "00010110001011101101101111100111100101110111011100000011001101010100000010010100111000011101100100010010" when "00010111010",
      "00010110010100011100001111010110101111001111011101101000000000011010000001100110010011001001101011000001" when "00010111011",
      "00010110011101001011000010001000111101100101101000111001100110010100110010011101001100110000000111000001" when "00010111100",
      "00010110100101111010000111111111100100000110110001110110001010111000101011010000100101011101101100001001" when "00010111101",
      "00010110100101111010000111111111100100000110110001110110001010111000101011010000100101011101101100001001" when "00010111110",
      "00010110101110101001100000111011110110001000001101110101111001111001100000010001001001001101010110110000" when "00010111111",
      "00010110110111011001001100111111000111000111110100110101100000110100000101001000001101010000001100100100" when "00011000000",
      "00010111000000001001001100001010101010101100000010100000111101000110110101001100111011110110100110010010" when "00011000001",
      "00010111001000111001011110011111110100100011110111011110010111011100001001111111011110000100011011000111" when "00011000010",
      "00010111010001101010000011111111111000100110111010011001001011101001000111100001110111100010110110011101" when "00011000011",
      "00010111010001101010000011111111111000100110111010011001001011101001000111100001110111100010110110011101" when "00011000100",
      "00010111011010011010111100101100001010110101011001001101011101100011000111001110110110101001010100111101" when "00011000101",
      "00010111100011001100001000100101111111011000001010010011011010101111001010010110110100111111011011100010" when "00011000110",
      "00010111101011111101100111101110101010100000101101101011001001001101011101110100001001000110100111101011" when "00011000111",
      "00010111110100101111011010000111100000101001001110001000100011000011111001110000011001110000011000111110" when "00011001000",
      "00010111111101100001011111110001110110010100100010011111011111001010000111111101011110100110100100000110" when "00011001001",
      "00010111111101100001011111110001110110010100100010011111011111001010000111111101011110100110100100000110" when "00011001010",
      "00011000000110010011111000101111000000001110001110110000000110111001111100101101111111111011111011101101" when "00011001011",
      "00011000001111000110100101000000010011001010100101010011011001000110101110100010011000111110100010110111" when "00011001100",
      "00011000010111111001100100100111000100000110101000000111111001111110011001101000111100111110001110001001" when "00011001101",
      "00011000100000101100110111100100101000001000001001111110110000010110111100111001000111101100110100111110" when "00011001110",
      "00011000100000101100110111100100101000001000001001111110110000010110111100111001000111101100110100111110" when "00011001111",
      "00011000101001100000011101111010010100011101101111101000110000001010111110011011110101101101111101110000" when "00011010000",
      "00011000110010010100010111101001011110011110110001000011110010001000000110111100111111111100101000101110" when "00011010001",
      "00011000111011001000100100110011011011101011011010101000011000110010000011001100000001000010101011000110" when "00011010010",
      "00011001000011111101000101011001100001101100101110010111100010111100111011111100000001011010110010101010" when "00011010011",
      "00011001001100110001111001011101000110010100100101001000101011100001110101011110101000111110110011001101" when "00011010100",
      "00011001001100110001111001011101000110010100100101001000101011100001110101011110101000111110110011001101" when "00011010101",
      "00011001010101100111000000111111011111011101101111110111110110110000000111111111000011011011001110101010" when "00011010110",
      "00011001011110011100011100000010000011001011111000110100001100111110100011001101111101101100001100011000" when "00011010111",
      "00011001100111010010001010100110000111101011100100101110100010111110110000011010001000101000010011000110" when "00011011000",
      "00011001110000001000001100101101000011010010010100001000001111110110000101111100011110011001100000101010" when "00011011001",
      "00011001111000111110100010011000001100011110100100100010010000011110100001001010000101011100111000010000" when "00011011010",
      "00011001111000111110100010011000001100011110100100100010010000011110100001001010000101011100111000010000" when "00011011011",
      "00011010000001110101001011101000111001110111110001101100011000110010011011001010010101011100100000010111" when "00011011100",
      "00011010001010101100001000100000100010001110010110110100110010100110001110011010110111110110111111000011" when "00011011101",
      "00011010010011100011011001000000011100011011101111110111101010010010100011010111011111110000011011110111" when "00011011110",
      "00011010011100011010111101001001111111100010011010101111001001010001111011001000000001111110111110101010" when "00011011111",
      "00011010011100011010111101001001111111100010011010101111001001010001111011001000000001111110111110101010" when "00011100000",
      "00011010100101010010110100111110100010101101111000100011011110010100110000000010110001001010111101010110" when "00011100001",
      "00011010101110001011000000011111011101010010101110111011010011101110100100011110100111010110000011011100" when "00011100010",
      "00011010110111000011011111101110000110101110101001001100010011011111011000111100111001101111101110011001" when "00011100011",
      "00011010111111111100010010101011110110101000011001101011111001011100000011011111110010101100110100101101" when "00011100100",
      "00011010111111111100010010101011110110101000011001101011111001011100000011011111110010101100110100101101" when "00011100101",
      "00011011001000110101011001011010000100101111111011000000010011011000100010101111011001000111110000110110" when "00011100110",
      "00011011010001101110110011111010001000111110010001010001101111010111000111111101000101100010001011000010" when "00011100111",
      "00011011011010101000100010001101011011010101101011011011110111111111010100000010001001011100011010110101" when "00011101000",
      "00011011100011100010100100010101010100000001100100011111011110111111100100000100011111011110110001000011" when "00011101001",
      "00011011101100011100111010010011001011010110100100110100010101111100101010111010011001000111001000100001" when "00011101010",
      "00011011101100011100111010010011001011010110100100110100010101111100101010111010011001000111001000100001" when "00011101011",
      "00011011110101010111100100001000011001110010100011011011010101010001110101110100001001111001100001000110" when "00011101100",
      "00011011111110010010100001110110010111111100100111010000110001100100011011000001001000010100000110001110" when "00011101101",
      "00011100000111001101110011011110011110100101001000011110111111001110010001110100000001000110111001101111" when "00011101110",
      "00011100010000001001011001000010000110100101110001110001000100100001110100011001001100001101110010001011" when "00011101111",
      "00011100010000001001011001000010000110100101110001110001000100100001110100011001001100001101110010001011" when "00011110000",
      "00011100011001000101010010100010101001000001100001100101111010001010101100100000110001001110010110100010" when "00011110001",
      "00011100100010000001100000000001011111000100101011100011011010001110001100101101010101100110100110011100" when "00011110010",
      "00011100101010111110000001100000000010000100111001101001111101101110011000100111101000010000010101100100" when "00011110011",
      "00011100110011111010110110111111101011100001001101101000001000110010111111100111000100100101010110100110" when "00011110100",
      "00011100110011111010110110111111101011100001001101101000001000110010111111100111000100100101010110100110" when "00011110101",
      "00011100111100111000000000100001110101000010000010001110100101011011001101101110111011001100101101111000" when "00011110110",
      "00011101000101110101011110000111111000011001001100100100001100111011010111101111101111101110110101011010" when "00011110111",
      "00011101001110110011001111110011001111100001111101011010100000001001100111101101001010000000001110110100" when "00011111000",
      "00011101010111110001010101100101010100100001000010100010001110011100110000011000010101000110100101010010" when "00011111001",
      "00011101010111110001010101100101010100100001000010100010001110011100110000011000010101000110100101010010" when "00011111010",
      "00011101100000101111101111011111100001100100101000000000001011100000001110100000010000110100101010000000" when "00011111011",
      "00011101101001101110011101100011010001000100011001100010010100000000011111101001110001011100110011000000" when "00011111100",
      "00011101110010101101011111110001111101100001100011110101000001010010110111010010001111001010101011111010" when "00011111101",
      "00011101110010101101011111110001111101100001100011110101000001010010110111010010001111001010101011111010" when "00011111110",
      "00011101111011101100110110001101000001100110110101111000101011111011111011010001011001011000101110000001" when "00011111111",
      "00011110000100101100100000110101111000001000100010010111011101010111110010000000000011001111110010010000" when "00100000000",
      "00011110001101101100011111101101111100000100100000111011010000100111001100111011001101010101111001110110" when "00100000001",
      "00011110010110101100110010110110101000100010001111100100000010000100111011001101001101100101011111010111" when "00100000010",
      "00011110010110101100110010110110101000100010001111100100000010000100111011001101001101100101011111010111" when "00100000011",
      "00011110011111101101011010010001011000110010110011111110001110100110010000111000100001000000011001100010" when "00100000100",
      "00011110101000101110010101111111101000010000111100111001100001101010001111110010001100010011110100011010" when "00100000101",
      "00011110110001101111100110000010110010100001000011011111110010111010100000001100110111010000111111100110" when "00100000110",
      "00011110111010110001001010011100010011010001001100101100010011000001001000000111100100011111001100100100" when "00100000111",
      "00011110111010110001001010011100010011010001001100101100010011000001001000000111100100011111001100100100" when "00100001000",
      "00011111000011110011000011001101100110011001001010100011000111110110110000100111001011000001110111001010" when "00100001001",
      "00011111001100110101010000011000000111111010011101101000111000001100001001110100001001011110110111011110" when "00100001010",
      "00011111010101110111110001111101010100000000010110011010100110110010011110101010001011000001001101101100" when "00100001011",
      "00011111010101110111110001111101010100000000010110011010100110110010011110101010001011000001001101101100" when "00100001100",
      "00011111011110111010100111111110100110111111110110100101111101000101101010011010100110001000011100111101" when "00100001101",
      "00011111100111111101110010011101011101010111110010100001100101011100000010110110111010110001100111111101" when "00100001110",
      "00011111110001000001010001011011010011110000110010100101110100111110101010101100100010010000000111011111" when "00100001111",
      "00011111111010000101000100111001100110111101010100100101100101001101100000101111011110101000000110110010" when "00100010000",
      "00011111111010000101000100111001100110111101010100100101100101001101100000101111011110101000000110110010" when "00100010001",
      "00100000000011001001001100111001110011111001101101000111011101010011000001000110100001101110000101100000" when "00100010010",
      "00100000001100001101101001011101010111101100001000111111001011001010001110011111111100111011111111001000" when "00100010011",
      "00100000010101010010011010100101101111100100101110100111001100011010111010101011010011011001010110000000" when "00100010100",
      "00100000010101010010011010100101101111100100101110100111001100011010111010101011010011011001010110000000" when "00100010101",
      "00100000011110010111100000010100011000111101011111011010100111001111000101101001111111000101101111101000" when "00100010110",
      "00100000100111011100111010101010110001011010011001001111010011000101001100011110000000010000000010101010" when "00100010111",
      "00100000110000100010101001101010010110101001010111110000010001100010100000110100000011101110100101001110" when "00100011000",
      "00100000111001101000101101010100100110100010010101111000010111001001000011111100010010001001101010011100" when "00100011001",
      "00100000111001101000101101010100100110100010010101111000010111001001000011111100010010001001101010011100" when "00100011010",
      "00100001000010101111000101101010111111000111001111001101000100010100011111111011001101111110101000000110" when "00100011011",
      "00100001001011110101110010101110111110100100000001011001101110100001011011010011001010010100010000001011" when "00100011100",
      "00100001010100111100110100100010000011001110101101101010111001100010100011111100110111101101011100111010" when "00100011101",
      "00100001010100111100110100100010000011001110101101101010111001100010100011111100110111101101011100111010" when "00100011110",
      "00100001011110000100001011000101101011100111011010001010000001000111001110111101100111000010100101001111" when "00100011111",
      "00100001100111001011110110011011010110011000010011011001010010110110101011111111110101010001000110110101" when "00100100000",
      "00100001110000010011110110100100100010010101101101101111111000100011101011101011010101001001101110101000" when "00100100001",
      "00100001111001011100001011100010101110011110000110110110010010111011111001010001011110010011101101000011" when "00100100010",
      "00100001111001011100001011100010101110011110000110110110010010111011111001010001011110010011101101000011" when "00100100011",
      "00100010000010100100110101010111011001111010000111000011000100110110101000111010001011000101110100000010" when "00100100100",
      "00100010001011101101110100000100000011111100100010110111101111000110011100010110100000111111100011100110" when "00100100101",
      "00100010010100110111000111101010001100000010011100011101111100110001000001010110100001011100101110011100" when "00100100110",
      "00100010010100110111000111101010001100000010011100011101111100110001000001010110100001011100101110011100" when "00100100111",
      "00100010011110000000110000001011010001110011000101000101000000010001001101011000010011010111101110100100" when "00100101000",
      "00100010100111001010101101101000110100111111111110011111100001000110011011011111111000011001000111000010" when "00100101001",
      "00100010110000010101000000000100010101100100111100100001011010010101010010000000010011110001111010100000" when "00100101010",
      "00100010110000010101000000000100010101100100111100100001011010010101010010000000010011110001111010100000" when "00100101011",
      "00100010111001011111100111011111010011101000000110011110001001111100110110011000001100010111111111010010" when "00100101100",
      "00100011000010101010100011111011001111011001111000100111010001000100010110111101100110110100100011010001" when "00100101101",
      "00100011001011110101110101011001101001010101000101101011000101000100110010101111011001110011011001110011" when "00100101110",
      "00100011001011110101110101011001101001010101000101101011000101000100110010101111011001110011011001110011" when "00100101111",
      "00100011010101000001011011111100000001111110111000010011110001110010001000011100010011001001101000100001" when "00100110000",
      "00100011011110001101010111100011111010000110110100100110101100100111110111001010101010100010110000001001" when "00100110001",
      "00100011100111011001101000010010110010100110111001100011111000111100011011100110110101010000011100010101" when "00100110010",
      "00100011100111011001101000010010110010100110111001100011111000111100011011100110110101010000011100010101" when "00100110011",
      "00100011110000100110001110001010001100100011100010100101111101011111010101111000110110000000110110111101" when "00100110100",
      "00100011111001110011001001001011101001001011101001000010001011000101100100111101111100100111001101011001" when "00100110101",
      "00100100000011000000011001011000101001111000100101101000110100101000000101011101110010101111101010000011" when "00100110110",
      "00100100000011000000011001011000101001111000100101101000110100101000000101011101110010101111101010000011" when "00100110111",
      "00100100001100001101111110110010110000001110010010000101111000011000000010101111001110001111111011011010" when "00100111000",
      "00100100010101011011111001011011011101111011001010100001111010101100101001111100101101001111000000000100" when "00100111001",
      "00100100011110101010001001010100010100111000001111000011010010001110001111110100111101111101011100010101" when "00100111010",
      "00100100100111111000101110011110110111001001000101001111100101100010011010110001000011010010111111001010" when "00100111011",
      "00100100100111111000101110011110110111001001000101001111100101100010011010110001000011010010111111001010" when "00100111100",
      "00100100110001000111101000111100100110111011111001101101011010011101000011110110000111000010011111100001" when "00100111101",
      "00100100111010010110111000101111000110101001100001100110010110111010000010010110011101011001001001001001" when "00100111110",
      "00100101000011100110011101110111111000110101011100001001010011100011010110010011000000101110011001101000" when "00100111111",
      "00100101000011100110011101110111111000110101011100001001010011100011010110010011000000101110011001101000" when "00101000000",
      "00100101001100110110011000011000100000001101110100001101000000000111100111011100000010001101100010101000" when "00101000001",
      "00100101010110000110101000010010011111101011100001110010111001100100101111001110010011011101011000001110" when "00101000010",
      "00100101010110000110101000010010011111101011100001110010111001100100101111001110010011011101011000001110" when "00101000011",
      "00100101011111010111001101100111011010010010001011101010010010001010100101001000000110100100110101110000" when "00101000100",
      "00100101101000101000001000011000110011010000001000110011101011011001100101110000001101101001010000011010" when "00101000101",
      "00100101110001111001011000101000001101111110100010000100100010000001001110001000000000001011011100101101" when "00101000110",
      "00100101110001111001011000101000001101111110100010000100100010000001001110001000000000001011011100101101" when "00101000111",
      "00100101111011001010111110010111001110000001010011101011001100000010000101100000111101000000110101010111" when "00101001000",
      "00100110000100011100111001100111010111000111001110110011001000110111110001001101100001010011110111000011" when "00101001001",
      "00100110001101101111001010011010001101001001111011001001100011101110001110100101000010000000111111001101" when "00101001010",
      "00100110001101101111001010011010001101001001111011001001100011101110001110100101000010000000111111001101" when "00101001011",
      "00100110010111000001110000110001010100001101111000100010001000000110110000110010011100010001010010111010" when "00101001100",
      "00100110100000010100101100101110010000100010100000011100001000110000100000100110001011000111100110011000" when "00101001101",
      "00100110101001100111111110010010100110100010000111100111111000111000011101100011111101010110110011111111" when "00101001110",
      "00100110101001100111111110010010100110100010000111100111111000111000011101100011111101010110110011111111" when "00101001111",
      "00100110110010111011100101011111111010110001111111101100010111110101000001000110100101101110010100010011" when "00101010000",
      "00100110111100001111100010010111110010000010011000101101001111010001000100110100110001111001011111101111" when "00101010001",
      "00100111000101100011110100111011110001001110100010110001000011111010101110100011111010000000011100001010" when "00101010010",
      "00100111000101100011110100111011110001001110100010110001000011111010101110100011111010000000011100001010" when "00101010011",
      "00100111001110111000011101001101011101011100101111100111111000111001100101100111010010101111100010100100" when "00101010100",
      "00100111011000001101011011001110011011111110010100010010000101110000110101101100110111110000010100100110" when "00101010101",
      "00100111100001100010101111000000010010001111101010100111011111010001000101001010100010110101111010010101" when "00101010110",
      "00100111100001100010101111000000010010001111101010100111011111010001000101001010100010110101111010010101" when "00101010111",
      "00100111101010111000011000100100100101111000010010111110110010111110000101000010010110110001001011000101" when "00101011000",
      "00100111110100001110010111111100111100101010110101110101010101101100100010100110101010010010010001110000" when "00101011001",
      "00100111110100001110010111111100111100101010110101110101010101101100100010100110101010010010010001110000" when "00101011010",
      "00100111111101100100101101001010111100100101000101010111000100111100000011001010111001010101100101111101" when "00101011011",
      "00101000000110111011011000010000001011101111111111000110111011010001010011110001001111011110110110100001" when "00101011100",
      "00101000010000010010011001001110010000011111101101100111010111110100110111101001011111011101111011101011" when "00101011101",
      "00101000010000010010011001001110010000011111101101100111010111110100110111101001011111011101111011101011" when "00101011110",
      "00101000011001101001110000000110110001010011101010000011011000111010100001011001110000101010111011010101" when "00101011111",
      "00101000100011000001011100111011010100110110011101110111101001110101100011101110010011111001111001110010" when "00101100000",
      "00101000101100011001011111101101100001111110000100011100000011111110000111110010101110000000100100111000" when "00101100001",
      "00101000101100011001011111101101100001111110000100011100000011111110000111110010101110000000100100111000" when "00101100010",
      "00101000110101110001111000011110111111101011101100101101100011001011111000011011110111101111100101110000" when "00101100011",
      "00101000111111001010100111010001010101001011111010111000001101101010010010001111110111111100111010011101" when "00101100100",
      "00101001001000100011101100000110001001110110101010000001101111001010101001111110110110110011110000111011" when "00101100101",
      "00101001001000100011101100000110001001110110101010000001101111001010101001111110110110110011110000111011" when "00101100110",
      "00101001010001111101000110111111000101001111001101110100000111111000011011100101110111010111001000101000" when "00101100111",
      "00101001011011010110110111111101101111000100010100001000101110110011110101011011100111100101010001101011" when "00101101000",
      "00101001011011010110110111111101101111000100010100001000101110110011110101011011100111100101010001101011" when "00101101001",
      "00101001100100110000111111000011101111010000000110110011100111110111010100001101101110111011001100000001" when "00101101010",
      "00101001101110001011011100010010101101111000001101001111001101101100000101011100001111111110000111010000" when "00101101011",
      "00101001110111100110001111101100010011001101101110001000001111010010000111001000110011010101001100100110" when "00101101100",
      "00101001110111100110001111101100010011001101101110001000001111010010000111001000110011010101001100100110" when "00101101101",
      "00101010000001000001011001010010000111101101010001001010000001011111111100110110101000100101101101111000" when "00101101110",
      "00101010001010011100111001000101110011111111000000101011000100011110110011000000110101110111101100110010" when "00101101111",
      "00101010001010011100111001000101110011111111000000101011000100011110110011000000110101110111101100110010" when "00101110000",
      "00101010010011111000101111001001000000110110101011011001111101000111001010110100101111101110001101010010" when "00101110001",
      "00101010011101010100111011011101010111010011100110001010100010100010101010000111001001011101010100000000" when "00101110010",
      "00101010100110110001011110000100100000100000101101100011011111110111001011100100011010000110110000011000" when "00101110011",
      "00101010100110110001011110000100100000100000101101100011011111110111001011100100011010000110110000011000" when "00101110100",
      "00101010110000001110010111000000000101110100100111101100001010000000001101000100110011101100101111011000" when "00101110101",
      "00101010111001101011100110010001110000110001100101111010101001111010011010111000100001111111011000011100" when "00101110110",
      "00101010111001101011100110010001110000110001100101111010101001111010011010111000100001111111011000011100" when "00101110111",
      "00101011000011001001001011111011001011000101100110100010011011000110010111101000110010110100010001011100" when "00101111000",
      "00101011001100100111000111111101111110101010010110100010111110100110100010010110001101011111101011010100" when "00101111001",
      "00101011010110000101011010011011110101100101010011010111000010011101011100100111010111110011011000110100" when "00101111010",
      "00101011010110000101011010011011110101100101010011010111000010011101011100100111010111110011011000110100" when "00101111011",
      "00101011011111100100000011010110011010000111101100100011111101110000010100100101110110011111100100000100" when "00101111100",
      "00101011101001000011000010101111010110101110100101101001100001010010110111010011011100111101010111011111" when "00101111101",
      "00101011101001000011000010101111010110101110100101101001100001010010110111010011011100111101010111011111" when "00101111110",
      "00101011110010100010011000101000010110000010110111110001111101000000110001001101011011110001010110000100" when "00101111111",
      "00101011111100000010000101000011000010111001010011100010011010001001100011111111110000011011101110111000" when "00110000000",
      "00101100000101100010001000000001001000010010100010101011101010010011011001110111000001111110101111111010" when "00110000001",
      "00101100000101100010001000000001001000010010100010101011101010010011011001110111000001111110101111111010" when "00110000010",
      "00101100001111000010100001100100010001011011001001111011001011011001011111101100110110000110000010000010" when "00110000011",
      "00101100011000100011010001101110001001101011101010101100100000101010110000110111100001010110010010111111" when "00110000100",
      "00101100011000100011010001101110001001101011101010101100100000101010110000110111100001010110010010111111" when "00110000101",
      "00101100100010000100011000100000011100101000100100111011000000101101100000010100000011001000101011110011" when "00110000110",
      "00101100101011100101110101111100110110000010011000110011111000101100101100001111000010111001110111100100" when "00110000111",
      "00101100110101000111101010000101000001110101101000101000100100110011101010100000000000101001011111111001" when "00110001000",
      "00101100110101000111101010000101000001110101101000101000100100110011101010100000000000101001011111111001" when "00110001001",
      "00101100111110101001110100111010101100001010111010100001011101111100111101011000111110010010110100000010" when "00110001010",
      "00101101001000001100010110011111100001010110111010010000111100111001000001011011110010110011000011101011" when "00110001011",
      "00101101001000001100010110011111100001010110111010010000111100111001000001011011110010110011000011101011" when "00110001100",
      "00101101010001101111001110110101001101111010011011000110110010110001100110010101111010100101100110100001" when "00110001101",
      "00101101011011010010011101111101011110100010011001100011110111001110100110010011010011100000010010110010" when "00110001110",
      "00101101011011010010011101111101011110100010011001100011110111001110100110010011010011100000010010110010" when "00110001111",
      "00101101100100110110000011111010000000000111111101001110001100000001010000001001100100110100100011011001" when "00110010000",
      "00101101101110011010000000101100011111110000011010100101010110011010011010001100111110010011000110001000" when "00110010001",
      "00101101110111111110010100010110101010101101010100110111001110010000110100110001111011110000111101001100" when "00110010010",
      "00101101110111111110010100010110101010101101010100110111001110010000110100110001111011110000111101001100" when "00110010011",
      "00101110000001100010111110111010001110011100011111110101000010111100010100101111010101011100110111011000" when "00110010100",
      "00101110001011001000000000011000111000101000000001101000110110001010101111100111011000011100000111000100" when "00110010101",
      "00101110001011001000000000011000111000101000000001101000110110001010101111100111011000011100000111000100" when "00110010110",
      "00101110010100101101011000110100010111000110010100101011001100110011100100001111001110001110000010100111" when "00110010111",
      "00101110011110010011001000001110010111111010001001011001010101101111001011111111111110100101100110001000" when "00110011000",
      "00101110011110010011001000001110010111111010001001011001010101101111001011111111111110100101100110001000" when "00110011001",
      "00101110100111111001001110101000101001010010101000001011100110110110110010001110110100001000111100111000" when "00110011010",
      "00101110110001011111101100000100111001101011010011001100010000010001110000011101000001100000111101111111" when "00110011011",
      "00101110110001011111101100000100111001101011010011001100010000010001110000011101000001100000111101111111" when "00110011100",
      "00101110111011000110100000100100110111101100001000001110100101110101101111100100110100011100111101111111" when "00110011101",
      "00101111000100101101101100001010010010001001100010100110011110111110001111011011101011110011111011001000" when "00110011110",
      "00101111001110010101001110110110111000000100011101000000001101000000110111010111100111000010111100110101" when "00110011111",
      "00101111001110010101001110110110111000000100011101000000001101000000110111010111100111000010111100110101" when "00110100000",
      "00101111010111111101001000101100011000101010010011011000101000000011010011111001100000011010100011000110" when "00110100001",
      "00101111100001100101011001101100100011010101000100110101110010011000000110110100010111100000111111101011" when "00110100010",
      "00101111100001100101011001101100100011010101000100110101110010011000000110110100010111100000111111101011" when "00110100011",
      "00101111101011001110000001111001000111101011010101011111110010100111010000011110011111110001010010010000" when "00110100100",
      "00101111110100110111000001010011110101100000010000011010000100100111111010010000001110010011110000000000" when "00110100101",
      "00101111110100110111000001010011110101100000010000011010000100100111111010010000001110010011110000000000" when "00110100110",
      "00101111111110100000010111111110011100110011101001011101000001010000001011101010000100100000101110100000" when "00110100111",
      "00110000001000001010000101111010101101110001111111001111111101000000010100110011010000010111001100100011" when "00110101000",
      "00110000001000001010000101111010101101110001111111001111111101000000010100110011010000010111001100100011" when "00110101001",
      "00110000010001110100001011001010011000110100011101000011011101101110011010011000110001111010000011000100" when "00110101010",
      "00110000011011011110100111101111001110100000111100101100000111010111110000101101000101100111011010110101" when "00110101011",
      "00110000100101001001011011101010111111101010001000011101011111111101010100100000011110011111011100000110" when "00110101100",
      "00110000100101001001011011101010111111101010001000011101011111111101010100100000011110011111011100000110" when "00110101101",
      "00110000101110110100100110111111011101001111011101000101101010110000010010000011000000011011101000011100" when "00110101110",
      "00110000111000100000001001101110011000011101001011101000111010110100001011111001101011110111010100010101" when "00110101111",
      "00110000111000100000001001101110011000011101001011101000111010110100001011111001101011110111010100010101" when "00110110000",
      "00110001000010001100000011111001100010101100011011011101111100111011110100101010000111000100101100010110" when "00110110001",
      "00110001001011111000010101100010101101100011001100001010011001000110001111111001101000001011000100100001" when "00110110010",
      "00110001001011111000010101100010101101100011001100001010011001000110001111111001101000001011000100100001" when "00110110011",
      "00110001010101100100111110101011101010110100010111011111101011100001010000010111010100011010001111011110" when "00110110100",
      "00110001011111010001111111010110001100011111110011011000010101010110101010100010110110100110010111101001" when "00110110101",
      "00110001011111010001111111010110001100011111110011011000010101010110101010100010110110100110010111101001" when "00110110110",
      "00110001101000111111010111100100000100110010010011110101100101001001110100011101010111001000100101111001" when "00110110111",
      "00110001110010101101000111010111000110000101101100111101010111001010101100101101000100010100000000001000" when "00110111000",
      "00110001110010101101000111010111000110000101101100111101010111001010101100101101000100010100000000001000" when "00110111001",
      "00110001111100011011001110110001000011000000110100111000101101100100000100011000011001110110010011110000" when "00110111010",
      "00110010000110001001101101110011101110010111100101110010100000101010001000111001110010100000110101101101" when "00110111011",
      "00110010000110001001101101110011101110010111100101110010100000101010001000111001110010100000110101101101" when "00110111100",
      "00110010001111111000100100100000111011001010111111110110100111001111001100001010000111000011000110011110" when "00110111101",
      "00110010011001100111110010111010011100101001001011010001010111000011101010111101010001111101100110011010" when "00110111110",
      "00110010011001100111110010111010011100101001001011010001010111000011101010111101010001111101100110011010" when "00110111111",
      "00110010100011010111011001000010000110001101011010001111011101100111010011001010000000101011100110110001" when "00111000000",
      "00110010101101000111010110111001101011100000001010111110010001010000101100010100000111111110110111101001" when "00111000001",
      "00110010101101000111010110111001101011100000001010111110010001010000101100010100000111111110110111101001" when "00111000010",
      "00110010110110110111101100100011000000010111001001101100011010110001000111001111011011110010101100101111" when "00111000011",
      "00110011000000101000011001111111111000110101010010101010110111011001111010010000010001011110001000010101" when "00111000100",
      "00110011000000101000011001111111111000110101010010101010110111011001111010010000010001011110001000010101" when "00111000101",
      "00110011001010011001011111010010001001001010110100001110010011101001010001011110010111110001001001110010" when "00111000110",
      "00110011010100001010111100011011100101110101010000110000111110100011111011111110110000111000111111000100" when "00111000111",
      "00110011010100001010111100011011100101110101010000110000111110100011111011111110110000111000111111000100" when "00111001000",
      "00110011011101111100110001011110000011011111100000110100110110000001100000001001111001101101010011100000" when "00111001001",
      "00110011100111101110111110011011010111000001110101000110001011110001000011000100000101001110001101110000" when "00111001010",
      "00110011100111101110111110011011010111000001110101000110001011110001000011000100000101001110001101110000" when "00111001011",
      "00110011110001100001100011010101010101100001111000011110100011011011110000001111101101001010101110001100" when "00111001100",
      "00110011111011010100100000001101110100010010110010001000001001101011010000110010110000001011110011010000" when "00111001101",
      "00110011111011010100100000001101110100010010110010001000001001101011010000110010110000001011110011010000" when "00111001110",
      "00110100000101000111110101000110101000110101000111100001100100011001100010001011001011100011000100101000" when "00111001111",
      "00110100001110111011100010000001101000110110111110100001111100001111111110110000110010000111111100111000" when "00111010000",
      "00110100001110111011100010000001101000110110111110100001111100001111111110110000110010000111111100111000" when "00111010001",
      "00110100011000101111100111000000101010010011111111011101011111011011101011100110010100001101010110110010" when "00111010010",
      "00110100100010100100000100000101100011010101010111001010011101111100100000011111011100010111000011010011" when "00111010011",
      "00110100100010100100000100000101100011010101010111001010011101111100100000011111011100010111000011010011" when "00111010100",
      "00110100101100011000111001010010001010010001111001000110011111010101000001000101010100011011000010100010" when "00111010101",
      "00110100110110001110000110101000010101101110000001011100010010000000111111001000010011110011101001010110" when "00111010110",
      "00110100110110001110000110101000010101101110000001011100010010000000111111001000010011110011101001010110" when "00111010111",
      "00110101000000000011101100001001111100011011110111001001110100011000011111110010100100111100110000011000" when "00111011000",
      "00110101001001111001101001111000110101011011001110000110110111100101011111010100111011110100101110010000" when "00111011001",
      "00110101001001111001101001111000110101011011001110000110110111100101011111010100111011110100101110010000" when "00111011010",
      "00110101010011101111111111110110110111111001101001001011111100010001110000001101100010101010100111011000" when "00111011011",
      "00110101011101100110101110000101111011010010011100011001101001010011010100001110101100110010011111010101" when "00111011100",
      "00110101011101100110101110000101111011010010011100011001101001010011010100001110101100110010011111010101" when "00111011101",
      "00110101100111011101110100100111110111001110101111000000011100011101001111110011001001110000001101111100" when "00111011110",
      "00110101110001010101010011011110100011100101011101101000110101011010111001010100111101010101000001000100" when "00111011111",
      "00110101110001010101010011011110100011100101011101101000110101011010111001010100111101010101000001000100" when "00111100000",
      "00110101111011001101001010101011111000011011011100011011111010111011101000000100001010110110010001001110" when "00111100001",
      "00110110000101000101011010010001101110000011011001001100011010010101000111100011001100111000100110001101" when "00111100010",
      "00110110000101000101011010010001101110000011011001001100011010010101000111100011001100111000100110001101" when "00111100011",
      "00110110001110111110000010010001111100111101111101100000000001100010010110010111111100110011100111110001" when "00111100100",
      "00110110011000110111000010101110011101111001110000111001010011100101011000101010011000111100101010110110" when "00111100101",
      "00110110011000110111000010101110011101111001110000111001010011100101011000101010011000111100101010110110" when "00111100110",
      "00110110100010110000011011101001001001110011011011000001110111110010001000010011100011111100001010001010" when "00111100111",
      "00110110101100101010001101000011111001110101100101110101000011101000001110101010100100011101111010000100" when "00111101000",
      "00110110101100101010001101000011111001110101100101110101000011101000001110101010100100011101111010000100" when "00111101001",
      "00110110110110100100010111000000100111011000111111101010111111100010010101001000011010011011100110001110" when "00111101010",
      "00110111000000011110111001100001001100000100011101100100000110100000111011100111001101011101100111110001" when "00111101011",
      "00110111000000011110111001100001001100000100011101100100000110100000111011100111001101011101100111110001" when "00111101100",
      "00110111001010011001110100100111100001101100111101010101000000110111000101101101101001000101000110000100" when "00111101101",
      "00110111001010011001110100100111100001101100111101010101000000110111000101101101101001000101000110000100" when "00111101110",
      "00110111010100010101001000010101100010010101100111110010111001111111010001000100001100101101101000010110" when "00111101111",
      "00110111011110010000110100101101001000001111110011000000010001011110101000111111001001100010001111111001" when "00111110000",
      "00110111011110010000110100101101001000001111110011000000010001011110101000111111001001100010001111111001" when "00111110001",
      "00110111101000001100111001110000001101111011000100011010000111011101001101010101111101101010010100010111" when "00111110010",
      "00110111110010001001010111100000101110000101010011000101100100011001000100001111010100000101100110100110" when "00111110011",
      "00110111110010001001010111100000101110000101010011000101100100011001000100001111010100000101100110100110" when "00111110100",
      "00110111111100000110001110000000100011101010101001111101111100011011001111110111101010110101001101111000" when "00111110101",
      "00111000000110000011011101010001101001110101101010000011001110010100100011100111111101010110100111111010" when "00111110110",
      "00111000000110000011011101010001101001110101101010000011001110010100100011100111111101010110100111111010" when "00111110111",
      "00111000010000000001000101010101111011111111001100101000111110001000110101010001110000101001110100110000" when "00111111000",
      "00111000011001111111000110001111010101101110100101100101101011101111001000110111000000101000101100110000" when "00111111001",
      "00111000011001111111000110001111010101101110100101100101101011101111001000110111000000101000101100110000" when "00111111010",
      "00111000100011111101011111111111110010111001100101100010100101001101010111100100010011100111011001010011" when "00111111011",
      "00111000101101111100010010101001001111100100011100001011110101010101110011110110100001011000111010111110" when "00111111100",
      "00111000101101111100010010101001001111100100011100001011110101010101110011110110100001011000111010111110" when "00111111101",
      "00111000110111111011011110001101101000000001111010100001001110001101001110100110100111010100001011011011" when "00111111110",
      "00111000110111111011011110001101101000000001111010100001001110001101001110100110100111010100001011011011" when "00111111111",
      "00111001000001111011000010101110111000110011010101000111010000000000000011001001010010100000111010110000" when "01000000000",
      "00111001001011111011000000001110111110101000100110011000101100001101010001100011011100110110001001110111" when "01000000001",
      "00111001001011111011000000001110111110101000100110011000101100001101010001100011011100110110001001110111" when "01000000010",
      "00111001010101111011010110101111110110100000010000111000100101001101110000101000010000111000111110000100" when "01000000011",
      "00111001011111111100000110010011011101100111100001100100101010011110100010101010000101000000000111001010" when "01000000100",
      "00111001011111111100000110010011011101100111100001100100101010011110100010101010000101000000000111001010" when "01000000101",
      "00111001101001111101001110111011110001011010010010001000010001010100111001111100011101110011000100111110" when "01000000110",
      "00111001110011111110110000101010101111100011001011001111101010100010111011111011001101010111010110100001" when "01000000111",
      "00111001110011111110110000101010101111100011001011001111101010100010111011111011001101010111010110100001" when "01000001000",
      "00111001111110000000101011100010010101111011100110111011110100110011010011100000001110010001000001111010" when "01000001001",
      "00111001111110000000101011100010010101111011100110111011110100110011010011100000001110010001000001111010" when "01000001010",
      "00111010001000000010111111100100100010101011110010110110101100000011000101001001001000010010001110001101" when "01000001011",
      "00111010010010000101101100110011010100001010110010100111110110000000011001000100100000111011011111010011" when "01000001100",
      "00111010010010000101101100110011010100001010110010100111110110000000011001000100100000111011011111010011" when "01000001101",
      "00111010011100001000110011010000101000111110100010001001101011110100110001110110110011010100001111110100" when "01000001110",
      "00111010100110001100010010111110011111111011110111111111000001000010000111011111001010010001110111111110" when "01000001111",
      "00111010100110001100010010111110011111111011110111111111000001000010000111011111001010010001110111111110" when "01000010000",
      "00111010110000010000001011111110111000000110100111101001000111111001000000111101111100101100011100100100" when "01000010001",
      "00111010111010010100011110010011110000110001100011111110010011001111101000010111110111001110000010111101" when "01000010010",
      "00111010111010010100011110010011110000110001100011111110010011001111101000010111110111001110000010111101" when "01000010011",
      "00111011000100011001001001111111001001011110100001100000110101111111110111001011010000001010111100000100" when "01000010100",
      "00111011000100011001001001111111001001011110100001100000110101111111110111001011010000001010111100000100" when "01000010101",
      "00111011001110011110001111000011000001111110011000110110100000010011111010100111111010010011000110010110" when "01000010110",
      "00111011011000100011101101100001011010010001001001000000011010101000010001110101001001111110010110110011" when "01000010111",
      "00111011011000100011101101100001011010010001001001000000011010101000010001110101001001111110010110110011" when "01000011000",
      "00111011100010101001100101011100010010100101111001110011011110101010001001001110000110000001011011100110" when "01000011001",
      "00111011101100101111110110110101101011011010111110010001001110011001011000111000101010010001010011011010" when "01000011010",
      "00111011101100101111110110110101101011011010111110010001001110011001011000111000101010010001010011011010" when "01000011011",
      "00111011110110110110100001101111100101011101110111000001001001010101001101011001010110001001011110010111" when "01000011100",
      "00111011110110110110100001101111100101011101110111000001001001010101001101011001010110001001011110010111" when "01000011101",
      "00111100000000111101100110001100000001101011010100101010011111111010100100100011011101011110111000000111" when "01000011110",
      "00111100001011000101000100001101000001001111011010001110100101011011101001100100010101010010011010000111" when "01000011111",
      "00111100001011000101000100001101000001001111011010001110100101011011101001100100010101010010011010000111" when "01000100000",
      "00111100010101001100111011110100100101100101011111100011100000010111011110000111000010000001100110101111" when "01000100001",
      "00111100011111010101001101000100110000011000010011101111011001011000111111101110000000101111111111011100" when "01000100010",
      "00111100011111010101001101000100110000011000010011101111011001011000111111101110000000101111111111011100" when "01000100011",
      "00111100101001011101110111111111100011100001111111100100001001000100111011000000100000111110100001100000" when "01000100100",
      "00111100101001011101110111111111100011100001111111100100001001000100111011000000100000111110100001100000" when "01000100101",
      "00111100110011100110111100100111000001001100000111111011100100011101100000001010101010001110110001001100" when "01000100110",
      "00111100111101110000011010111101001011101111110000010100001000100011101110010000110110010011011011101011" when "01000100111",
      "00111100111101110000011010111101001011101111110000010100001000100011101110010000110110010011011011101011" when "01000101000",
      "00111101000111111010010011000100000101110101011101001110000100111101001100111001100000011110010100011010" when "01000101001",
      "00111101010010000100100100111101110010010101010110101001000101100110001101110011001010100011010111111100" when "01000101010",
      "00111101010010000100100100111101110010010101010110101001000101100110001101110011001010100011010111111100" when "01000101011",
      "00111101011100001111010000101100010100010111001010100010011011110111010010000000100010110111111110100100" when "01000101100",
      "00111101011100001111010000101100010100010111001010100010011011110111010010000000100010110111111110100100" when "01000101101",
      "00111101100110011010010110010001101111010010001111010011100111000101110000011000101010011011111110011010" when "01000101110",
      "00111101110000100101110101110000000110101101100110010001011100100110111101001101111000100110000100111100" when "01000101111",
      "00111101110000100101110101110000000110101101100110010001011100100110111101001101111000100110000100111100" when "01000110000",
      "00111101111010110001101111001001011110011111111110001011101111011101010100110100100010001110001111011110" when "01000110001",
      "00111101111010110001101111001001011110011111111110001011101111011101010100110100100010001110001111011110" when "01000110010",
      "00111110000100111110000010011111111010101111110101101101010111110111001101000111111101010101101100101001" when "01000110011",
      "00111110001111001010101111110101011111110011011101111100111010100110110100010011111000000100100110001101" when "01000110100",
      "00111110001111001010101111110101011111110011011101111100111010100110110100010011111000000100100110001101" when "01000110101",
      "00111110011001010111110111001100010010010000111100111101110000011011000100101111100010110000010001010000" when "01000110110",
      "00111110100011100101011000100110010110111110010000010001101101100000111000100000100001001010001001010101" when "01000110111",
      "00111110100011100101011000100110010110111110010000010001101101100000111000100000100001001010001001010101" when "01000111000",
      "00111110101101110011010100000101110011000001001111011011001001010100101001000011110110100110001010000010" when "01000111001",
      "00111110101101110011010100000101110011000001001111011011001001010100101001000011110110100110001010000010" when "01000111010",
      "00111110111000000001101001101100101011101111101110011111100110101011101001100110001100000111011101011010" when "01000111011",
      "00111111000010010000011001011101000110101111100000101010111100011101001100111101100111100011011010111100" when "01000111100",
      "00111111000010010000011001011101000110101111100000101010111100011101001100111101100111100011011010111100" when "01000111101",
      "00111111001100011111100011011001001001110110011010110010111110110011001010000011001101111100110000000101" when "01000111110",
      "00111111001100011111100011011001001001110110011010110010111110110011001010000011001101111100110000000101" when "01000111111",
      "00111111010110101111000111100010111011001010010101111011101001001001110011110101111100001011011101101001" when "01001000000",
      "00111111100000111111000101111100100001000001010001111011101001000110111100011100111101101001111110011110" when "01001000001",
      "00111111100000111111000101111100100001000001010001111011101001000110111100011100111101101001111110011110" when "01001000010",
      "00111111101011001111011110101000000010000001011000000001101010001111111100101100110011000100010101000101" when "01001000011",
      "00111111101011001111011110101000000010000001011000000001101010001111111100101100110011000100010101000101" when "01001000100",
      "00111111110101100000010001100111100101000000111101011010000011000110111100000000010010011100010110100110" when "01001000101",
      "00111111111111110001011110111101010001000110100101110101000011010110110110100101001110101101000111100000" when "01001000110",
      "00111111111111110001011110111101010001000110100101110101000011010110110110100101001110101101000111100000" when "01001000111",
      "01000000001010000011000110101011001101101001000110001101100011010110100010001011100111100001011110101000" when "01001001000",
      "01000000010100010101001000110011100010001111100111010000010101001010110011110110100010111101101000001111" when "01001001001",
      "01000000010100010101001000110011100010001111100111010000010101001010110011110110100010111101101000001111" when "01001001010",
      "01000000011110100111100101011000010110110001101000000011110111001111101011011110100001011010110110011010" when "01001001011",
      "01000000011110100111100101011000010110110001101000000011110111001111101011011110100001011010110110011010" when "01001001100",
      "01000000101000111010011100011011110011010111000000110000101000110000101100000110011001110111111111110110" when "01001001101",
      "01000000110011001101101110000000000000011000000101001001111111111000101010010110011000111001010111000111" when "01001001110",
      "01000000110011001101101110000000000000011000000101001001111111111000101010010110011000111001010111000111" when "01001001111",
      "01000000111101100001011010000111000110011101100111010111100010000000111100100011011000010000100011001011" when "01001010000",
      "01000000111101100001011010000111000110011101100111010111100010000000111100100011011000010000100011001011" when "01001010001",
      "01000001000111110101100000110011001110100000111010011110111110001000011010011100101111111001111000110100" when "01001010010",
      "01000001010010001010000010000110100001101011110101001110101001011010011100101110111011011001110001100111" when "01001010011",
      "01000001010010001010000010000110100001101011110101001110101001011010011100101110111011011001110001100111" when "01001010100",
      "01000001011100011110111110000011001001011000110100101000011110001110001110111110011001011010110000110010" when "01001010101",
      "01000001011100011110111110000011001001011000110100101000011110001110001110111110011001011010110000110010" when "01001010110",
      "01000001100110110100010100101011001111010010111110101101011101100110101000110100100101001110001011111000" when "01001010111",
      "01000001110001001010000110000000111101010110000101001001110011011011000101101110110101001110100100010100" when "01001011000",
      "01000001110001001010000110000000111101010110000101001001110011011011000101101110110101001110100100010100" when "01001011001",
      "01000001111011100000010010000110011101101110101000000001011101010001110100110111000101001110010000010010" when "01001011010",
      "01000001111011100000010010000110011101101110101000000001011101010001110100110111000101001110010000010010" when "01001011011",
      "01000010000101110110111000111101111010111001111000011101010100010011111101000101111111100111101010011000" when "01001011100",
      "01000010010000001101111010101001011111100101111011011000111010000011110011100111010111000000110111111010" when "01001011101",
      "01000010010000001101111010101001011111100101111011011000111010000011110011100111010111000000110111111010" when "01001011110",
      "01000010011010100101010111001011010110110001101100010000101000011110000101110011010000110100001001101010" when "01001011111",
      "01000010011010100101010111001011010110110001101100010000101000011110000101110011010000110100001001101010" when "01001100000",
      "01000010100100111101001110100101101011101100111111110000100101001110011001101001000011000100001110111111" when "01001100001",
      "01000010101111010101100000111010101001111000100110100011111000011111101010010100011011000000010011011111" when "01001100010",
      "01000010101111010101100000111010101001111000100110100011111000011111101010010100011011000000010011011111" when "01001100011",
      "01000010111001101110001110001100011101000110010000000100100111010001001001000001000111110010100000000010" when "01001100100",
      "01000010111001101110001110001100011101000110010000000100100111010001001001000001000111110010100000000010" when "01001100101",
      "01000011000100000111010110011101010001011000101101001100010001011000101100011110011101010111010001001000" when "01001100110",
      "01000011000100000111010110011101010001011000101101001100010001011000101100011110011101010111010001001000" when "01001100111",
      "01000011001110100000111001101111010011000011110011000100110011011010111100010001101110111110001011101100" when "01001101000",
      "01000011011000111010111000000100101110101100011101111010001100100010000111010100111111101000110101000010" when "01001101001",
      "01000011011000111010111000000100101110101100011101111010001100100010000111010100111111101000110101000010" when "01001101010",
      "01000011100011010101010001011111110001001000110011101100101000011100010111011110111001010100100110110000" when "01001101011",
      "01000011100011010101010001011111110001001000110011101100101000011100010111011110111001010100100110110000" when "01001101100",
      "01000011101101110000000110000010100111100000000111000011001101101010010110110000100001101011111010101000" when "01001101101",
      "01000011111000001011010101101111011111001010111001111111010000000110111101000110111101110100111111001110" when "01001101110",
      "01000011111000001011010101101111011111001010111001111111010000000110111101000110111101110100111111001110" when "01001101111",
      "01000100000010100111000000101000100101110011000000110000001000010001000000010000000101001011110011010010" when "01001110000",
      "01000100000010100111000000101000100101110011000000110000001000010001000000010000000101001011110011010010" when "01001110001",
      "01000100001101000011000110110000001001010011100100100111101111000000000001100100100111011100011100100100" when "01001110010",
      "01000100010111011111101000001000010111111001000110101111011110001100111000101101000001111111000111001100" when "01001110011",
      "01000100010111011111101000001000010111111001000110101111011110001100111000101101000001111111000111001100" when "01001110100",
      "01000100100001111100100100110011100000000001100010111101110110010111011011111010101111011010010010111101" when "01001110101",
      "01000100100001111100100100110011100000000001100010111101110110010111011011111010101111011010010010111101" when "01001110110",
      "01000100101100011001111100110011110000011100010010101100101001010010001010000100011111011110010111010001" when "01001110111",
      "01000100101100011001111100110011110000011100010010101100101001010010001010000100011111011110010111010001" when "01001111000",
      "01000100110110110111110000001011011000001010001111101111101001111100111100011010011111011011000000010100" when "01001111001",
      "01000101000001010101111110111100100110011101110111001100000001111000001001001101101010101111010100111110" when "01001111010",
      "01000101000001010101111110111100100110011101110111001100000001111000001001001101101010101111010100111110" when "01001111011",
      "01000101001011110100101001001001101010111011001100010000001011111001000010101101000010111100010001110000" when "01001111100",
      "01000101001011110100101001001001101010111011001100010000001011111001000010101101000010111100010001110000" when "01001111101",
      "01000101010110010011101110110100110101010111111011001100010100101001000000100100101010100010111011011000" when "01001111110",
      "01000101100000110011010000000000010101111011011100001011100000111000100100110010110100001001001100000111" when "01001111111",
      "01000101100000110011010000000000010101111011011100001011100000111000100100110010110100001001001100000111" when "01010000000",
      "01000101101011010011001100101110011100111110110110001101011001101111101111010010100010110100000010010100" when "01010000001",
      "01000101101011010011001100101110011100111110110110001101011001101111101111010010100010110100000010010100" when "01010000010",
      "01000101110101110011100101000001011011001101000010000000011111000100110110100101011101010010111101001010" when "01010000011",
      "01000101110101110011100101000001011011001101000010000000011111000100110110100101011101010010111101001010" when "01010000100",
      "01000110000000010100011000111011100001100010101100111101000000000011011110010010110001110001101010011000" when "01010000101",
      "01000110001010110101101000011111000001001110011100000000011010001100100110111110011100111111111011010101" when "01010000110",
      "01000110001010110101101000011111000001001110011100000000011010001100100110111110011100111111111011010101" when "01010000111",
      "01000110010101010111010011101110001011110000101110101001011110111001110101101000110101010000101000010110" when "01010001000",
      "01000110010101010111010011101110001011110000101110101001011110111001110101101000110101010000101000010110" when "01010001001",
      "01000110011111111001011010101011010010111100000001110100111111101100110011110110000000101101110101000000" when "01010001010",
      "01000110011111111001011010101011010010111100000001110100111111101100110011110110000000101101110101000000" when "01010001011",
      "01000110101010011011111101011000101000110100110010111011000001010100101100001011011110111100111111111010" when "01010001100",
      "01000110110100111110111011111000011111110001100010101100110101110011001001100011001000000001111101010110" when "01010001101",
      "01000110110100111110111011111000011111110001100010101100110101110011001001100011001000000001111101010110" when "01010001110",
      "01000110111111100010010110001101001010011010111000010011011101101010100010100011110111101101101101101111" when "01010001111",
      "01000110111111100010010110001101001010011010111000010011011101101010100010100011110111101101101101101111" when "01010010000",
      "01000111001010000110001100011000111011101011100100001110110000011110111101000010101010100110010100100100" when "01010010001",
      "01000111001010000110001100011000111011101011100100001110110000011110111101000010101010100110010100100100" when "01010010010",
      "01000111010100101010011110011110000110110000100011010101001100110011111000100001011100101011011001110010" when "01010010011",
      "01000111011111001111001100011110111111001001000001110100001111110000010001010101111101111110001110010100" when "01010010100",
      "01000111011111001111001100011110111111001001000001110100001111110000010001010101111101111110001110010100" when "01010010101",
      "01000111101001110100010110011101111000100110011110010001010100010010110000110111010010011010000111100101" when "01010010110",
      "01000111101001110100010110011101111000100110011110010001010100010010110000110111010010011010000111100101" when "01010010111",
      "01000111110100011001111100011101000111001100101100101011011010100000000010000110101110101000110100000000" when "01010011000",
      "01000111110100011001111100011101000111001100101100101011011010100000000010000110101110101000110100000000" when "01010011001",
      "01000111111110111111111110011110111111010001111001011101010110110101000100111111111100001100000101000101" when "01010011010",
      "01001000001001100110011100100101110101011110101100100000101001100111011101010011100100101001101000011010" when "01010011011",
      "01001000001001100110011100100101110101011110101100100000101001100111011101010011100100101001101000011010" when "01010011100",
      "01001000010100001101010110110011111110101110001100010000111110111101011101001000110101110101110100110000" when "01010011101",
      "01001000010100001101010110110011111110101110001100010000111110111101011101001000110101110101110100110000" when "01010011110",
      "01001000011110110100101101001011110000001110000000110000010111001000001101111100000000011100010101011100" when "01010011111",
      "01001000011110110100101101001011110000001110000000110000010111001000001101111100000000011100010101011100" when "01010100000",
      "01001000101001011100011111101111011111011110010110101011110111101001111101101010011111110010011000101000" when "01010100001",
      "01001000110100000100101110100001100010010010000010100001000101010010011000111001000100101011010110001111" when "01010100010",
      "01001000110100000100101110100001100010010010000010100001000101010010011000111001000100101011010110001111" when "01010100011",
      "01001000111110101101011001100100001110101110100011100100000110111011011101011101000110101101110111111000" when "01010100100",
      "01001000111110101101011001100100001110101110100011100100000110111011011101011101000110101101110111111000" when "01010100101",
      "01001001001001010110100000111001111011001100000111000110010001110000110100001111100111111100010111000100" when "01010100110",
      "01001001001001010110100000111001111011001100000111000110010001110000110100001111100111111100010111000100" when "01010100111",
      "01001001010100000000000100100100111110010101101011011101011110101100000011101111011101111111001001010010" when "01010101000",
      "01001001011110101010000100100111101111001001000011001100001001010000001111110111011010111000110110010001" when "01010101001",
      "01001001011110101010000100100111101111001001000011001100001001010000001111110111011010111000110110010001" when "01010101010",
      "01001001101001010100100001000100100100110110111000001001111000001110111110101101110110011101101100000010" when "01010101011",
      "01001001101001010100100001000100100100110110111000001001111000001110111110101101110110011101101100000010" when "01010101100",
      "01001001110011111111011001111101110111000010101110101100110000000001011100110101000000000101001100111000" when "01010101101",
      "01001001110011111111011001111101110111000010101110101100110000000001011100110101000000000101001100111000" when "01010101110",
      "01001001111110101010101111010101111101100011001000110011001110111111111110100101101000010010110010011100" when "01010101111",
      "01001001111110101010101111010101111101100011001000110011001110111111111110100101101000010010110010011100" when "01010110000",
      "01001010001001010110100001001111010000100001101001001110110100000010011111100001011010010101001001100011" when "01010110001",
      "01001010010100000010101111101100001000011010110110101111001111010100100011001111000111010111010101000110" when "01010110010",
      "01001010010100000010101111101100001000011010110110101111001111010100100011001111000111010111010101000110" when "01010110011",
      "01001010011110101111011010101110111101111110011111001110011101100111011110111000010001001000011001111101" when "01010110100",
      "01001010011110101111011010101110111101111110011111001110011101100111011110111000010001001000011001111101" when "01010110101",
      "01001010101001011100100010011010001010001111011010111101001110001101010101000110101111010001100010010000" when "01010110110",
      "01001010101001011100100010011010001010001111011010111101001110001101010101000110101111010001100010010000" when "01010110111",
      "01001010110100001010000110110000000110100011101111110000010011100111010001101000011011000110000011100010" when "01010111000",
      "01001010111110111000000111110011001100100100110100001110011111010010010100101000000000100111100111111000" when "01010111001",
      "01001010111110111000000111110011001100100100110100001110011111010010010100101000000000100111100111111000" when "01010111010",
      "01001011001001100110100101100101110110001111010010111111001000011101000001010011101010011010010010111110" when "01010111011",
      "01001011001001100110100101100101110110001111010010111111001000011101000001010011101010011010010010111110" when "01010111100",
      "01001011010100010101100000001010011101110011001101111001011110010001000110010101010111110011010100100001" when "01010111101",
      "01001011010100010101100000001010011101110011001101111001011110010001000110010101010111110011010100100001" when "01010111110",
      "01001011011111000100110111100011011101110100000001010100100101011011111001101100101011100010110010101000" when "01010111111",
      "01001011011111000100110111100011011101110100000001010100100101011011111001101100101011100010110010101000" when "01011000000",
      "01001011101001110100101011110011010001001000100111011000000001100000100101000110100011101110000011110110" when "01011000001",
      "01001011110100100100111100111100010010111011011011001101001001111111000010111110010011100000100110010000" when "01011000010",
      "01001011110100100100111100111100010010111011011011001101001001111111000010111110010011100000100110010000" when "01011000011",
      "01001011111111010101101011000000111110101010011100010001001011011010101111100001100100011101000111001010" when "01011000100",
      "01001011111111010101101011000000111110101010011100010001001011011010101111100001100100011101000111001010" when "01011000101",
      "01001100001010000110110110000011110000000111010001100111110100101100010100100001110111101011010100100010" when "01011000110",
      "01001100001010000110110110000011110000000111010001100111110100101100010100100001110111101011010100100010" when "01011000111",
      "01001100010100111000011110000111000011010111001101001110110000101001011001101111011000011010001111000010" when "01011001000",
      "01001100010100111000011110000111000011010111001101001110110000101001011001101111011000011010001111000010" when "01011001001",
      "01001100011111101010100011001101010100110011001111010001101100001101100111001011010000101101110000111000" when "01011001010",
      "01001100011111101010100011001101010100110011001111010001101100001101100111001011010000101101110000111000" when "01011001011",
      "01001100101010011101000101011001000001001000001001011111001001010000001001110011010111101011101011000101" when "01011001100",
      "01001100110101010000000100101100100101010110100010011101111110010001001110011101111110010010010011101100" when "01011001101",
      "01001100110101010000000100101100100101010110100010011101111110010001001110011101111110010010010011101100" when "01011001110",
      "01001101000000000011100001001010011110110010111001000011100011001010101010010001110101101110001011100101" when "01011001111",
      "01001101000000000011100001001010011110110010111001000011100011001010101010010001110101101110001011100101" when "01011010000",
      "01001101001010110111011010110101001011000101100111101010101011001111001010111110000111111101110101100100" when "01011010001",
      "01001101001010110111011010110101001011000101100111101010101011001111001010111110000111111101110101100100" when "01011010010",
      "01001101010101101011110001101111001000001011000111101011001100100011101101001101100001111000101111111001" when "01011010011",
      "01001101010101101011110001101111001000001011000111101011001100100011101101001101100001111000101111111001" when "01011010100",
      "01001101100000100000100101111010110100010011110100110010010100111110011010001001011101111010000111100010" when "01011010101",
      "01001101100000100000100101111010110100010011110100110010010100111110011010001001011101111010000111100010" when "01011010110",
      "01001101101011010101110111011010101110000100010000011011101100110110110000111100010111011111000111101010" when "01011010111",
      "01001101110110001011100110010001010100010101000101001011000111110010100100011101110010110101011000111110" when "01011011000",
      "01001101110110001011100110010001010100010101000101001011000111110010100100011101110010110101011000111110" when "01011011001",
      "01001110000001000001110010100001000110010011001010000111000011011011011000101111110001111110101001101110" when "01011011010",
      "01001110000001000001110010100001000110010011001010000111000011011011011000101111110001111110101001101110" when "01011011011",
      "01001110001011111000011100001100100011011111100110010011110100101000001111010010101000101101101000100010" when "01011011100",
      "01001110001011111000011100001100100011011111100110010011110100101000001111010010101000101101101000100010" when "01011011101",
      "01001110010110101111100011010110001011101111110100001111100011000111010100110011100100110011100001011110" when "01011011110",
      "01001110010110101111100011010110001011101111110100001111100011000111010100110011100100110011100001011110" when "01011011111",
      "01001110100001100111001000000000011111001101100101001110110011110011100110011010101111011000110100111111" when "01011100000",
      "01001110100001100111001000000000011111001101100101001110110011110011100110011010101111011000110100111111" when "01011100001",
      "01001110101100011111001010001101111110010111000100111010000010000010000111111110101000001101101011000001" when "01011100010",
      "01001110110111010111101010000001001001111110111100101011100111110011001000100101100011111001011011001010" when "01011100011",
      "01001110110111010111101010000001001001111110111100101011100111110011001000100101100011111001011011001010" when "01011100100",
      "01001111000010010000100111011100100011001100010111001110110101010010110110000001101011110101011100010100" when "01011100101",
      "01001111000010010000100111011100100011001100010111001110110101010010110110000001101011110101011100010100" when "01011100110",
      "01001111001101001010000010100010101011011011000011111111010111110110000011011001000001101000001100111001" when "01011100111",
      "01001111001101001010000010100010101011011011000011111111010111110110000011011001000001101000001100111001" when "01011101000",
      "01001111011000000011111011010110000100011011011010101001110000011110101010110001011001000010111000110111" when "01011101001",
      "01001111011000000011111011010110000100011011011010101001110000011110101010110001011001000010111000110111" when "01011101010",
      "01001111100010111110010001111001010000010010011110101100011010010100010101011111011011010001101000101000" when "01011101011",
      "01001111100010111110010001111001010000010010011110101100011010010100010101011111011011010001101000101000" when "01011101100",
      "01001111101101111001000110001110110001011010000010111001100000111101011010000000110100111100000100001000" when "01011101101",
      "01001111101101111001000110001110110001011010000010111001100000111101011010000000110100111100000100001000" when "01011101110",
      "01001111111000110100011000011001001010100000101100111001100111000100100010010011101110011111000110010000" when "01011101111",
      "01010000000011110000001000011010111110101001111000101110111101010111010001001000011100110000100000110010" when "01011110000",
      "01010000000011110000001000011010111110101001111000101110111101010111010001001000011100110000100000110010" when "01011110001",
      "01010000001110101100010110010110110001001101111100011001101010001010000000010111010101111111011001010011" when "01011110010",
      "01010000001110101100010110010110110001001101111100011001101010001010000000010111010101111111011001010011" when "01011110011",
      "01010000011001101001000010001111000101111010001011011100100001101101110110010010000111000001001110011100" when "01011110100",
      "01010000011001101001000010001111000101111010001011011100100001101101110110010010000111000001001110011100" when "01011110101",
      "01010000100100100110001100000110100000110000111010100010101111100100110011010111000101010001001001000101" when "01011110110",
      "01010000100100100110001100000110100000110000111010100010101111100100110011010111000101010001001001000101" when "01011110111",
      "01010000101111100011110011111111100110001001100011000110010001000000111101111101001100110101010001000101" when "01011111000",
      "01010000101111100011110011111111100110001001100011000110010001000000111101111101001100110101010001000101" when "01011111001",
      "01010000111010100001111001111100111010110000100110110111000000111011010101000000111111000100011011001101" when "01011111010",
      "01010000111010100001111001111100111010110000100110110111000000111011010101000000111111000100011011001101" when "01011111011",
      "01010001000101100000011110000001000011100111110011100010110101001110110110101101101110000100111100000110" when "01011111100",
      "01010001000101100000011110000001000011100111110011100010110101001110110110101101101110000100111100000110" when "01011111101",
      "01010001010000011111100000001110100110000110000110011110001110000100101011110010001100110011011110101110" when "01011111110",
      "01010001011011011111000000101000000111110111110000001101110110111110001100000101111010101111010110100010" when "01011111111",
      "01010001011011011111000000101000000111110111110000001101110110111110001100000101111010101111010110100010" when "01100000000",
      "01010001100110011110111111010000001110111110011000010000111010001001110100111010010101110000100100110100" when "01100000001",
      "01010001100110011110111111010000001110111110011000010000111010001001110100111010010101110000100100110100" when "01100000010",
      "01010001110001011111011100001001100001110001000000101100000110001111101101001100000101001100010101101111" when "01100000011",
      "01010001110001011111011100001001100001110001000000101100000110001111101101001100000101001100010101101111" when "01100000100",
      "01010001111100100000010111010110100110111100001001110101100110100010111000000001001111000110101101011111" when "01100000101",
      "01010001111100100000010111010110100110111100001001110101100110100010111000000001001111000110101101011111" when "01100000110",
      "01010010000111100001110000111010000101100001110110000001101110000100011001011100111100100101111101001100" when "01100000111",
      "01010010000111100001110000111010000101100001110110000001101110000100011001011100111100100101111101001100" when "01100001000",
      "01010010010010100011101000110110100100111001101101010000010101100101010101101100011100001101111000010110" when "01100001001",
      "01010010010010100011101000110110100100111001101101010000010101100101010101101100011100001101111000010110" when "01100001010",
      "01010010011101100101111111001110101100110001000000111011001100110100110110101111010010111001100110101010" when "01100001011",
      "01010010011101100101111111001110101100110001000000111011001100110100110110101111010010111001100110101010" when "01100001100",
      "01010010101000101000110100000101000101001010101111100100111111000111101000011011100100011010000110100101" when "01100001101",
      "01010010101000101000110100000101000101001010101111100100111111000111101000011011100100011010000110100101" when "01100001110",
      "01010010110011101100000111011100010110011111101000101001001011100101111110111110101101010001100001010000" when "01100001111",
      "01010010110011101100000111011100010110011111101000101001001011100101111110111110101101010001100001010000" when "01100010000",
      "01010010111110101111111001010111001001011110010000001100110001001101111111111101110001011000111110101110" when "01100010001",
      "01010011001001110100001001111000000111001011000010101111101110110111001001111010100100111010111000010110" when "01100010010",
      "01010011001001110100001001111000000111001011000010101111101110110111001001111010100100111010111000010110" when "01100010011",
      "01010011010100111000111001000001111001000000011000111111010111100100111010100111110001010001000001011010" when "01100010100",
      "01010011010100111000111001000001111001000000011000111111010111100100111010100111110001010001000001011010" when "01100010101",
      "01010011011111111110000110110111001000101110101011101001011011010101111000011011101110000111011111000011" when "01100010110",
      "01010011011111111110000110110111001000101110101011101001011011010101111000011011101110000111011111000011" when "01100010111",
      "01010011101011000011110011011010100000011100010111010000000100011101000110111001010111100101111011001110" when "01100011000",
      "01010011101011000011110011011010100000011100010111010000000100011101000110111001010111100101111011001110" when "01100011001",
      "01010011110110001001111110101110101010100101111111111110101001110011010011001110110110110100011011011100" when "01100011010",
      "01010011110110001001111110101110101010100101111111111110101001110011010011001110110110110100011011011100" when "01100011011",
      "01010100000001010000101000110110010001111110010101011111010110001101101001010011111010011010110100010000" when "01100011100",
      "01010100000001010000101000110110010001111110010101011111010110001101101001010011111010011010110100010000" when "01100011101",
      "01010100001100010111110001110100000001101110010110110001100101001000000101111101100000111101001111101101" when "01100011110",
      "01010100001100010111110001110100000001101110010110110001100101001000000101111101100000111101001111101101" when "01100011111",
      "01010100010111011111011001101010100101010101010110000001010100110000111111101001011000111011001011110101" when "01100100000",
      "01010100010111011111011001101010100101010101010110000001010100110000111111101001011000111011001011110101" when "01100100001",
      "01010100100010100111100000011100101000101000111100011111001110000100000010110010011000111010110010110100" when "01100100010",
      "01010100100010100111100000011100101000101000111100011111001110000100000010110010011000111010110010110100" when "01100100011",
      "01010100101101110000000110001100110111110101001110011001100010100010100011001110101111110110111011101111" when "01100100100",
      "01010100101101110000000110001100110111110101001110011001100010100010100011001110101111110110111011101111" when "01100100101",
      "01010100111000111001001010111101111111011100101110110110000000010111001000101010101000111110011011001110" when "01100100110",
      "01010100111000111001001010111101111111011100101110110110000000010111001000101010101000111110011011001110" when "01100100111",
      "01010101000100000010101110110010101100011000100011101100011100110011000000000100011010011100110101000010" when "01100101000",
      "01010101000100000010101110110010101100011000100011101100011100110011000000000100011010011100110101000010" when "01100101001",
      "01010101001111001100110001101101101011111000011001100010010101010011000000100100010000100101010001101110" when "01100101010",
      "01010101001111001100110001101101101011111000011001100010010101010011000000100100010000100101010001101110" when "01100101011",
      "01010101011010010111010011110001101011100010100111100111000111011010110110011111000010110100011111110101" when "01100101100",
      "01010101011010010111010011110001101011100010100111100111000111011010110110011111000010110100011111110101" when "01100101101",
      "01010101100101100010010101000001011001010100010011110001011111110100101011101011011100011101110011100110" when "01100101110",
      "01010101100101100010010101000001011001010100010011110001011111110100101011101011011100011101110011100110" when "01100101111",
      "01010101110000101101110101011111100011100001010110011101100000100011101000101001100000111101111000001100" when "01100110000",
      "01010101111011111001110101001110111000110100011110101011011110110111101110010111010100000011101110100101" when "01100110001",
      "01010101111011111001110101001110111000110100011110101011011110110111101110010111010100000011101110100101" when "01100110010",
      "01010110000111000110010100010010001000001111010101111111111000110001101101001001010001001011010110110110" when "01100110011",
      "01010110000111000110010100010010001000001111010101111111111000110001101101001001010001001011010110110110" when "01100110100",
      "01010110010010010011010010101100000001001010100100100100000010100101100001011010100100001100110001101110" when "01100110101",
      "01010110010010010011010010101100000001001010100100100100000010100101100001011010100100001100110001101110" when "01100110110",
      "01010110011101100000110000011111010011010101110101000111101100101010000011101001000000001100110110011100" when "01100110111",
      "01010110011101100000110000011111010011010101110101000111101100101010000011101001000000001100110110011100" when "01100111000",
      "01010110101000101110101101101110101110110111111001000011100001100100111101010000100000010011000001111111" when "01100111001",
      "01010110101000101110101101101110101110110111111001000011100001100100111101010000100000010011000001111111" when "01100111010",
      "01010110110011111101001010011101000100001110101100011100011101000001011000111100110011001111010111111010" when "01100111011",
      "01010110110011111101001010011101000100001110101100011100011101000001011000111100110011001111010111111010" when "01100111100",
      "01010110111111001100000110101101000100001111011010000111111011100000101001001011101100111111001000001000" when "01100111101",
      "01010110111111001100000110101101000100001111011010000111111011100000101001001011101100111111001000001000" when "01100111110",
      "01010111001010011011100010100001100000000110011111110001000011010011100100011111111010100100000110000000" when "01100111111",
      "01010111001010011011100010100001100000000110011111110001000011010011100100011111111010100100000110000000" when "01101000000",
      "01010111010101101011011101111101001001010111110001111110100110101011111011101011011100110100010001110110" when "01101000001",
      "01010111010101101011011101111101001001010111110001111110100110101011111011101011011100110100010001110110" when "01101000010",
      "01010111100000111011111001000010110001111110100000011001111111110100110010100001011110101101000001110010" when "01101000011",
      "01010111100000111011111001000010110001111110100000011001111111110100110010100001011110101101000001110010" when "01101000100",
      "01010111101100001100110011110101001100001101011001110111000110100001001000101001110100010111111011101100" when "01101000101",
      "01010111101100001100110011110101001100001101011001110111000110100001001000101001110100010111111011101100" when "01101000110",
      "01010111110111011110001110010111001010101110110000011101000000000000000100011100010001111001101100100101" when "01101000111",
      "01010111110111011110001110010111001010101110110000011101000000000000000100011100010001111001101100100101" when "01101001000",
      "01011000000010110000001000101011100000100100011101101111101001000101110110110111110011111101100100100011" when "01101001001",
      "01011000000010110000001000101011100000100100011101101111101001000101110110110111110011111101100100100011" when "01101001010",
      "01011000001110000010100010110101000001001000000110111010011010111001010011111000101010100100110110100101" when "01101001011",
      "01011000001110000010100010110101000001001000000110111010011010111001010011111000101010100100110110100101" when "01101001100",
      "01011000011001010101011100110110100000001011000000111011101010010100111111100001110110111011100011010010" when "01101001101",
      "01011000011001010101011100110110100000001011000000111011101010010100111111100001110110111011100011010010" when "01101001110",
      "01011000100100101000110110110010110001110110010100110001000010101011110101000000111001111100001110011100" when "01101001111",
      "01011000100100101000110110110010110001110110010100110001000010101011110101000000111001111100001110011100" when "01101010000",
      "01011000101111111100110000101100101010101011000011100100111011100000110001100111001010001111111111111101" when "01101010001",
      "01011000101111111100110000101100101010101011000011100100111011100000110001100111001010001111111111111101" when "01101010010",
      "01011000111011010001001010100110111111100010001010111100101010000001010010001010001110100000000010011000" when "01101010011",
      "01011000111011010001001010100110111111100010001010111100101010000001010010001010001110100000000010011000" when "01101010100",
      "01011001000110100110000100100100100101101100101001000111101110010010010110110100101100100110101110010110" when "01101010101",
      "01011001000110100110000100100100100101101100101001000111101110010010010110110100101100100110101110010110" when "01101010110",
      "01011001010001111011011110101000010010110011100001001111111100100000000101101010000001000100001100011010" when "01101010111",
      "01011001010001111011011110101000010010110011100001001111111100100000000101101010000001000100001100011010" when "01101011000",
      "01011001011101010001011000110100111100110111111111101010100010011111101001011011100010110111101110000000" when "01101011001",
      "01011001011101010001011000110100111100110111111111101010100010011111101001011011100010110111101110000000" when "01101011010",
      "01011001101000100111110011001101011010010011011110001010001001110011101111001001111001110010001010100101" when "01101011011",
      "01011001101000100111110011001101011010010011011110001010001001110011101111001001111001110010001010100101" when "01101011100",
      "01011001110011111110101101110100100001110111101000010001110110100011101001101100011110101001110111111100" when "01101011101",
      "01011001110011111110101101110100100001110111101000010001110110100011101001101100011110101001110111111100" when "01101011110",
      "01011001111111010110001000101101001010101110011111101001000011010101000111111001100000011010111010110111" when "01101011111",
      "01011001111111010110001000101101001010101110011111101001000011010101000111111001100000011010111010110111" when "01101100000",
      "01011010001010101110000011111010001100011010100000010000011010011001001110101011011101011101000000000110" when "01101100001",
      "01011010001010101110000011111010001100011010100000010000011010011001001110101011011101011101000000000110" when "01101100010",
      "01011010010110000110011111011110011110110110100100110111101100011100101101100100101000011111110100001100" when "01101100011",
      "01011010010110000110011111011110011110110110100100110111101100011100101101100100101000011111110100001100" when "01101100100",
      "01011010100001011111011011011100111010010110001011010100100101001100001001010111101011011101100011011100" when "01101100101",
      "01011010100001011111011011011100111010010110001011010100100101001100001001010111101011011101100011011100" when "01101100110",
      "01011010101100111000110111111000010111100101011000111010011101111100011101100011101001010111011001101000" when "01101100111",
      "01011010101100111000110111111000010111100101011000111010011101111100011101100011101001010111011001101000" when "01101101000",
      "01011010111000010010110100110011101111101000111110110011001110101000011010011011100100101000000110101000" when "01101101001",
      "01011010111000010010110100110011101111101000111110110011001110101000011010011011100100101000000110101000" when "01101101010",
      "01011011000011101101010010010001111011111110011110011000111101010011101010111101001000010011101111000000" when "01101101011",
      "01011011000011101101010010010001111011111110011110011000111101010011101010111101001000010011101111000000" when "01101101100",
      "01011011001111001000010000010101110110011100001101110000101100100100010010100111000010101000110110101000" when "01101101101",
      "01011011001111001000010000010101110110011100001101110000101100100100010010100111000010101000110110101000" when "01101101110",
      "01011011011010100011101111000010011001010001011100000110001001000011011000101111000101110101111100100110" when "01101101111",
      "01011011011010100011101111000010011001010001011100000110001001000011011000101111000101110101111100100110" when "01101110000",
      "01011011100101111111101110011010011111000110010110001000010110010101111100001000100010110110000110100011" when "01101110001",
      "01011011100101111111101110011010011111000110010110001000010110010101111100001000100010110110000110100011" when "01101110010",
      "01011011100101111111101110011010011111000110010110001000010110010101111100001000100010110110000110100011" when "01101110011",
      "01011011110001011100001110100001000010111100001010100111011011011110101110111110101000011001100111001000" when "01101110100",
      "01011011110001011100001110100001000010111100001010100111011011011110101110111110101000011001100111001000" when "01101110101",
      "01011011111100111001001111011001000000001101001110110011001111011010100000011011100001100011000010100011" when "01101110110",
      "01011011111100111001001111011001000000001101001110110011001111011010100000011011100001100011000010100011" when "01101110111",
      "01011100001000010110110001000101010010101101000010111011000101100111011110101010111000101000001110011100" when "01101111000",
      "01011100001000010110110001000101010010101101000010111011000101100111011110101010111000101000001110011100" when "01101111001",
      "01011100010011110100110011101000110110101000010110101110011011001001100001011111101001010001110001110011" when "01101111010",
      "01011100010011110100110011101000110110101000010110101110011011001001100001011111101001010001110001110011" when "01101111011",
      "01011100011111010011010111000110101000100101001101111110100100011100010010111111001100100100100101011000" when "01101111100",
      "01011100011111010011010111000110101000100101001101111110100100011100010010111111001100100100100101011000" when "01101111101",
      "01011100101010110010011011100001100101100011000101000001011100000100110001010000100111101001011100100000" when "01101111110",
      "01011100101010110010011011100001100101100011000101000001011100000100110001010000100111101001011100100000" when "01101111111",
      "01011100110110010010000000111100101010111010110101010101010010110011101001101100111111011001100011000110" when "01110000000",
      "01011100110110010010000000111100101010111010110101010101010010110011101001101100111111011001100011000110" when "01110000001",
      "01011101000001110010000111011010110110011110111010000101100001001010010011101110001100000101100101011000" when "01110000010",
      "01011101000001110010000111011010110110011110111010000101100001001010010011101110001100000101100101011000" when "01110000011",
      "01011101001101010010101110111111000110011011010100110000011010110011110110011011111110101100000000100011" when "01110000100",
      "01011101001101010010101110111111000110011011010100110000011010110011110110011011111110101100000000100011" when "01110000101",
      "01011101011000110011110111101100011001010101110001101110000100000100001010011011100000010100011001101100" when "01110000110",
      "01011101011000110011110111101100011001010101110001101110000100000100001010011011100000010100011001101100" when "01110000111",
      "01011101100100010101100001100101101110001101101100111000001001101110101110001011101010111101111010011000" when "01110001000",
      "01011101100100010101100001100101101110001101101100111000001001101110101110001011101010111101111010011000" when "01110001001",
      "01011101101111110111101100101110000100011100010110010010111011100111001001100001010010110001010111001010" when "01110001010",
      "01011101101111110111101100101110000100011100010110010010111011100111001001100001010010110001010111001010" when "01110001011",
      "01011101111011011010011001001000011011110100110110110111001001111101100010000000010001001001000111110100" when "01110001100",
      "01011101111011011010011001001000011011110100110110110111001001111101100010000000010001001001000111110100" when "01110001101",
      "01011110000110111101100110110111110100100100010100111101000110001000100111111011011111110110001111010010" when "01110001110",
      "01011110000110111101100110110111110100100100010100111101000110001000100111111011011111110110001111010010" when "01110001111",
      "01011110010010100001010101111111001111010001111001001000100110110000001001010011110010101000011111001100" when "01110010000",
      "01011110010010100001010101111111001111010001111001001000100110110000001001010011110010101000011111001100" when "01110010001",
      "01011110010010100001010101111111001111010001111001001000100110110000001001010011110010101000011111001100" when "01110010010",
      "01011110011110000101100110100001101100111110110010110110001111101001011101111110100010111011110000001110" when "01110010011",
      "01011110011110000101100110100001101100111110110010110110001111101001011101111110100010111011110000001110" when "01110010100",
      "01011110101001101010011000100010001111000110011101001001011101111001000101101111101011011110001010100010" when "01110010101",
      "01011110101001101010011000100010001111000110011101001001011101111001000101101111101011011110001010100010" when "01110010110",
      "01011110110101001111101100000011110111011110100011011011111000001011010111010111000001111110000101000110" when "01110010111",
      "01011110110101001111101100000011110111011110100011011011111000001011010111010111000001111110000101000110" when "01110011000",
      "01011111000000110101100001001001101000010111000110001101100011110111000100111000010100101100000011010010" when "01110011001",
      "01011111000000110101100001001001101000010111000110001101100011110111000100111000010100101100000011010010" when "01110011010",
      "01011111001100011011110111110110100100011010011111110110011110111100011111111101110000110010001111000011" when "01110011011",
      "01011111001100011011110111110110100100011010011111110110011110111100011111111101110000110010001111000011" when "01110011100",
      "01011111011000000010110000001101101110101101101001011000111111010011101110100000011110100111111011001110" when "01110011101",
      "01011111011000000010110000001101101110101101101001011000111111010011101110100000011110100111111011001110" when "01110011110",
      "01011111100011101010001010010010001010101111111111010101010111011101000101111111010010110100110000010111" when "01110011111",
      "01011111100011101010001010010010001010101111111111010101010111011101000101111111010010110100110000010111" when "01110100000",
      "01011111101111010010000110000110111100011011100110011110100001000110101001111011101111000011110111101110" when "01110100001",
      "01011111101111010010000110000110111100011011100110011110100001000110101001111011101111000011110111101110" when "01110100010",
      "01011111111010111010100011101111001000000101010000101111101101111001101111110110110101001100101100010010" when "01110100011",
      "01011111111010111010100011101111001000000101010000101111101101111001101111110110110101001100101100010010" when "01110100100",
      "01011111111010111010100011101111001000000101010000101111101101111001101111110110110101001100101100010010" when "01110100101",
      "01100000000110100011100011001101110010011100100010000011011110100011110001001011000011001101110011000011" when "01110100110",
      "01100000000110100011100011001101110010011100100010000011011110100011110001001011000011001101110011000011" when "01110100111",
      "01100000010010001101000100100110000000101011110101001011100000101101011001100110101111011000010111010100" when "01110101000",
      "01100000010010001101000100100110000000101011110101001011100000101101011001100110101111011000010111010100" when "01110101001",
      "01100000011101110111000111111010111000011000100000101001110011110011100110110010101011010001011100001010" when "01110101010",
      "01100000011101110111000111111010111000011000100000101001110011110011100110110010101011010001011100001010" when "01110101011",
      "01100000101001100001101101001111011111100010111011101010110101010101110011111010110010010100010010010100" when "01110101100",
      "01100000101001100001101101001111011111100010111011101010110101010101110011111010110010010100010010010100" when "01110101101",
      "01100000110101001100110100100110111100100110100011000000110100101100110010011011110110100000110101010110" when "01110101110",
      "01100000110101001100110100100110111100100110100011000000110100101100110010011011110110100000110101010110" when "01110101111",
      "01100001000000111000011110000100010110011001111110000000001110111101110111000111111100110110000010010100" when "01110110000",
      "01100001000000111000011110000100010110011001111110000000001110111101110111000111111100110110000010010100" when "01110110001",
      "01100001001100100100101001101010110100001111000011011101010010111110001001000100101011011101000111100100" when "01110110010",
      "01100001001100100100101001101010110100001111000011011101010010111110001001000100101011011101000111100100" when "01110110011",
      "01100001011000010001010111011101011101110010111110101010101101111001100110011001101110111100010011101011" when "01110110100",
      "01100001011000010001010111011101011101110010111110101010101101111001100110011001101110111100010011101011" when "01110110101",
      "01100001011000010001010111011101011101110010111110101010101101111001100110011001101110111100010011101011" when "01110110110",
      "01100001100011111110100111011111011011001110010100011001100000110001111000111100010011000010000010101101" when "01110110111",
      "01100001100011111110100111011111011011001110010100011001100000110001111000111100010011000010000010101101" when "01110111000",
      "01100001101111101100011001110011110101000101000111111001111111001000111011011011110110011001100111110000" when "01110111001",
      "01100001101111101100011001110011110101000101000111111001111111001000111011011011110110011001100111110000" when "01110111010",
      "01100001111011011010101110011101110100010110111111111101110111001011010110001111100010011101000100000110" when "01110111011",
      "01100001111011011010101110011101110100010110111111111101110111001011010110001111100010011101000100000110" when "01110111100",
      "01100010000111001001100101100000100010011111001011111011100011101111000001000000000111011011010010011101" when "01110111101",
      "01100010000111001001100101100000100010011111001011111011100011101111000001000000000111011011010010011101" when "01110111110",
      "01100010010010111000111110111111001001010100101000110010101000011001111101001001101100001011101001110010" when "01110111111",
      "01100010010010111000111110111111001001010100101000110010101000011001111101001001101100001011101001110010" when "01111000000",
      "01100010011110101000111010111100110011001010000110010001011000000110000011110010001000100111000101100100" when "01111000001",
      "01100010011110101000111010111100110011001010000110010001011000000110000011110010001000100111000101100100" when "01111000010",
      "01100010101010011001011001011100101010101110001011111011100110010110000111110101000010011010011010000000" when "01111000011",
      "01100010101010011001011001011100101010101110001011111011100110010110000111110101000010011010011010000000" when "01111000100",
      "01100010101010011001011001011100101010101110001011111011100110010110000111110101000010011010011010000000" when "01111000101",
      "01100010110110001010011010100001111011001011011110010010100011110000110100001100011111011100011111010000" when "01111000110",
      "01100010110110001010011010100001111011001011011110010010100011110000110100001100011111011100011111010000" when "01111000111",
      "01100011000001111011111110001111110000001000100011111110000101110110010100000110110111100101101011011100" when "01111001000",
      "01100011000001111011111110001111110000001000100011111110000101110110010100000110110111100101101011011100" when "01111001001",
      "01100011001101101110000100101001010101101000001010110110111010100101011010100101000011010100011111010101" when "01111001010",
      "01100011001101101110000100101001010101101000001010110110111010100101011010100101000011010100011111010101" when "01111001011",
      "01100011011001100000101101110001111000001001001101010010001000000101000100101010010100110111001100101101" when "01111001100",
      "01100011011001100000101101110001111000001001001101010010001000000101000100101010010100110111001100101101" when "01111001101",
      "01100011100101010011111001101100100100100110110111001101111000100111011000110111011000111011101100000000" when "01111001110",
      "01100011100101010011111001101100100100100110110111001101111000100111011000110111011000111011101100000000" when "01111001111",
      "01100011100101010011111001101100100100100110110111001101111000100111011000110111011000111011101100000000" when "01111010000",
      "01100011110001000111101000011100101000011000101011011111010011011011001100111100101010110000100000111100" when "01111010001",
      "01100011110001000111101000011100101000011000101011011111010011011011001100111100101010110000100000111100" when "01111010010",
      "01100011111100111011111010000101010001010010101001000001100010100001100010000101010110001110000111111010" when "01111010011",
      "01100011111100111011111010000101010001010010101001000001100010100001100010000101010110001110000111111010" when "01111010100",
      "01100100001000110000101110101001101101100101010000000110000101111100001110010100010011101111111011010111" when "01111010101",
      "01100100001000110000101110101001101101100101010000000110000101111100001110010100010011101111111011010111" when "01111010110",
      "01100100010100100110000110001101001011111101100111100110010100101011010001000110011100111110000011010100" when "01111010111",
      "01100100010100100110000110001101001011111101100111100110010100101011010001000110011100111110000011010100" when "01111011000",
      "01100100100000011100000000110010111011100101100010010110001011101110010111101010110000001101011010011100" when "01111011001",
      "01100100100000011100000000110010111011100101100010010110001011101110010111101010110000001101011010011100" when "01111011010",
      "01100100101100010010011110011110001100000011100100011000001011100000011100111111110100110000110101100010" when "01111011011",
      "01100100101100010010011110011110001100000011100100011000001011100000011100111111110100110000110101100010" when "01111011100",
      "01100100101100010010011110011110001100000011100100011000001011100000011100111111110100110000110101100010" when "01111011101",
      "01100100111000001001011111010010001101011011001000010010100100000010111000001000110011011111101010111000" when "01111011110",
      "01100100111000001001011111010010001101011011001000010010100100000010111000001000110011011111101010111000" when "01111011111",
      "01100101000100000001000011010010010000001100100100100101110000001110010010101111111111111010000110111000" when "01111100000",
      "01100101000100000001000011010010010000001100100100100101110000001110010010101111111111111010000110111000" when "01111100001",
      "01100101001111111001001010100001100101010101010001000100000000011111001000110100111110010110110100101110" when "01111100010",
      "01100101001111111001001010100001100101010101010001000100000000011111001000110100111110010110110100101110" when "01111100011",
      "01100101011011110001110101000011011110001111101100001010010101010011111001101101101101101110110001010100" when "01111100100",
      "01100101011011110001110101000011011110001111101100001010010101010011111001101101101101101110110001010100" when "01111100101",
      "01100101100111101011000010111011001100110011100000011010101001110011011001101110111110110001110010010001" when "01111100110",
      "01100101100111101011000010111011001100110011100000011010101001110011011001101110111110110001110010010001" when "01111100111",
      "01100101100111101011000010111011001100110011100000011010101001110011011001101110111110110001110010010001" when "01111101000",
      "01100101110011100100110100001100000011010101101001110111001110110001011010111111010010011000001111100100" when "01111101001",
      "01100101110011100100110100001100000011010101101001110111001110110001011010111111010010011000001111100100" when "01111101010",
      "01100101111111011111001000111001010100101000011011011111010110101000001011001001110011101011000100011000" when "01111101011",
      "01100101111111011111001000111001010100101000011011011111010110101000001011001001110011101011000100011000" when "01111101100",
      "01100110001011011010000001000110010011111011100100101101010010011101001011011011001100000100010010011111" when "01111101101",
      "01100110001011011010000001000110010011111011100100101101010010011101001011011011001100000100010010011111" when "01111101110",
      "01100110010111010101011100110110010100111100010110110101100000101000001111001001100110111111101110001000" when "01111101111",
      "01100110010111010101011100110110010100111100010110110101100000101000001111001001100110111111101110001000" when "01111110000",
      "01100110010111010101011100110110010100111100010110110101100000101000001111001001100110111111101110001000" when "01111110001",
      "01100110100011010001011100001100101011110101101010100111001101010011010101000011100010111110101010110001" when "01111110010",
      "01100110100011010001011100001100101011110101101010100111001101010011010101000011100010111110101010110001" when "01111110011",
      "01100110101111001101111111001100101101010000000101101110000101001010010110011101100110001100100001011101" when "01111110100",
      "01100110101111001101111111001100101101010000000101101110000101001010010110011101100110001100100001011101" when "01111110101",
      "01100110111011001011000101111001101110010010000000010101011010110001101111010111010111100111010000110010" when "01111110110",
      "01100110111011001011000101111001101110010010000000010101011010110001101111010111010111100111010000110010" when "01111110111",
      "01100111000111001000110000010111000100011111101010101100011110111011001001110001111011111001000000101000" when "01111111000",
      "01100111000111001000110000010111000100011111101010101100011110111011001001110001111011111001000000101000" when "01111111001",
      "01100111000111001000110000010111000100011111101010101100011110111011001001110001111011111001000000101000" when "01111111010",
      "01100111010011000110111110101000000101111011010010101100001100001111011110010111100111111010011111000011" when "01111111011",
      "01100111010011000110111110101000000101111011010010101100001100001111011110010111100111111010011111000011" when "01111111100",
      "01100111011111000101110000110000001001000101001001011110000110100101100011111101000011001101011001111110" when "01111111101",
      "01100111011111000101110000110000001001000101001001011110000110100101100011111101000011001101011001111110" when "01111111110",
      "01100111101011000101000110110010100100111011101001000100101110011101001111001110010011101110010001001110" when "01111111111",
      "10110110010100100011011111011010111010111110011011001111011101000100110000001110100011001000011011010010" when "10000000000",
      "10110110011010100011100000111010111100011110011100001011011101111001100100000101010110111010000101110101" when "10000000001",
      "10110110100000100011101011011011001111111111000010010000101011010000111001011101100110011111101010110000" when "10000000010",
      "10110110100000100011101011011011001111111111000010010000101011010000111001011101100110011111101010110000" when "10000000011",
      "10110110100110100011111110111100010000100010011011011000010000111101110110110001010111000001110101111010" when "10000000100",
      "10110110101100100100011011011110011001001100101111001110011011111000101000000010101010100100100101100000" when "10000000101",
      "10110110110010100101000001000010000101000011111111011101110101111000000011111100100111111010101111011101" when "10000000110",
      "10110110111000100101101111100111101111010000000111111011000011000001001100011110010111110111000000111100" when "10000000111",
      "10110110111110100110100111001111110010111010111110110000000000001100110111010111000000110101001011100100" when "10000001000",
      "10110111000100100111100111111010101011010000010100100111100011000011101010011011101001010110101011111000" when "10000001001",
      "10110111001010101000110001101000110011011101110100111000111011010000011000000010101001100110001100011011" when "10000001010",
      "10110111010000101010000100011010100110110011000101110011010101001001000111110001010100100110000011001001" when "10000001011",
      "10110111010000101010000100011010100110110011000101110011010101001001000111110001010100100110000011001001" when "10000001100",
      "10110111010110101011100000010000100000100001101000101001011101101111010111101011000010010110001010001011" when "10000001101",
      "10110111011100101101000101001010111011111100111001111101001000000111000010010011000100111110100111010110" when "10000001110",
      "10110111100010101110110011001010010100011010010001101010110100000100110101110100010100100101011001101011" when "10000001111",
      "10110111101000110000101010001111000101010001000011010101010110010100001000100011111111000111000001011100" when "10000010000",
      "10110111101110110010101010011001101001111010011110010001100001110100010111010110101011110011110001010000" when "10000010001",
      "10110111110100110100110011101010011101110001101101110001110010101110011010000001000100010101110011111100" when "10000010010",
      "10110111111010110111000110000001111100010011111001010001111010100001111010011111011000011111010110111100" when "10000010011",
      "10110111111010110111000110000001111100010011111001010001111010100001111010011111011000011111010110111100" when "10000010100",
      "10111000000000111001100001100000100001000000000100100010101101101010111011000001010100110011111011010100" when "10000010101",
      "10111000000110111100000110000110100111010111001111110101110010011111110111111001101000001100010010110000" when "10000010110",
      "10111000001100111110110011110100101010111100011000001001010001101000010001010010111000011010001001110000" when "10000010111",
      "10111000010011000001101010101011000111010100010111010011100111101100001001101101001010001110111000000010" when "10000011000",
      "10111000011001000100101010101010011000000110000100001111011000011100100101101010000110100000001011000110" when "10000011001",
      "10111000011111000111110011110010111000111010010011000111000011010101011001001111001010110110000000001101" when "10000011010",
      "10111000100101001011000110000101000101011011110101100000111001011000010000000111111010010110110001100010" when "10000011011",
      "10111000100101001011000110000101000101011011110101100000111001011000010000000111111010010110110001100010" when "10000011100",
      "10111000101011001110100001100001011001010111011010101010110100100001011100110100001000101001111011100111" when "10000011101",
      "10111000110001010010000110001000010000011011101111100110010000010110011011110000000000000101010111100100" when "10000011110",
      "10111000110111010101110011111010000110011001011111010100000100001110010111000110001010101111111100011100" when "10000011111",
      "10111000111101011001101010110111010111000011010011000000011110110100110111111110001101010010110001001101" when "10000100000",
      "10111001000011011101101011000000011110001101110010001111000011000111010001111011101001111011111000010010" when "10000100001",
      "10111001001001100001110100010101110111101111100011000110100110101100010101100100001010010111101010001100" when "10000100010",
      "10111001001111100110000110110111111111100001001010011101010001100110110111000101010111100010110100000101" when "10000100011",
      "10111001001111100110000110110111111111100001001010011101010001100110110111000101010111100010110100000101" when "10000100100",
      "10111001010101101010100010100111010001011101001100000100011111100011010101110101001111001101000110011110" when "10000100101",
      "10111001011011101111000111100100001001100000001010110101000010100000110001101001110000010101010110000011" when "10000100110",
      "10111001100001110011110101101111000011101000101000111011000110110100111011000111000001010001101000111000" when "10000100111",
      "10111001100111111000101101001000011011110111001000000010011000101100001011100100111100011011001011101100" when "10000101000",
      "10111001101101111101101101110000101110001110001001100010001011000101010010001111111010110011111011011010" when "10000101001",
      "10111001110100000010110111101000010110110010001110101001100000001001000011001001111110110101010010110100" when "10000101010",
      "10111001111010001000001010101111110001101001111000101011010010111110010101010100001100101010101001110010" when "10000101011",
      "10111001111010001000001010101111110001101001111000101011010010111110010101010100001100101010101001110010" when "10000101100",
      "10111010000000001101100111000111011010111101101001001010100010111010011101001010001001101000010001010110" when "10000101101",
      "10111010000110010011001100101111101110111000000010000110100000001110010000011011100111110111111001000010" when "10000101110",
      "10111010001100011000111011101001001001100101100110000110111010010000000000110010110000010111010111101000" when "10000101111",
      "10111010010010011110110011110100000111010100111000101000001111000010011010010111001010000011101110001100" when "10000110000",
      "10111010011000100100110101010001000100010110011110000111111100011000110011100000101010100011101111100100" when "10000110001",
      "10111010011110101011000000000000011100111100111100010000110010011000111011001110101010011001000110010110" when "10000110010",
      "10111010011110101011000000000000011100111100111100010000110010011000111011001110101010011001000110010110" when "10000110011",
      "10111010100100110001010100000010101101011100111010000111000111011010010011011011000101001101100011110000" when "10000110100",
      "10111010101010110111110001011000010010001101000000010101001101100011100100100010011100111011111010100010" when "10000110101",
      "10111010110000111110011000000001100111100101111001010111101001100101110111111100100101111001001110110000" when "10000110110",
      "10111010110111000101000111111111001010000010010001101001101011010110100110100011110001100011011100001000" when "10000110111",
      "10111010111101001100000001010001010101111110110111110001100111100111101001001010011101010110000110011111" when "10000111000",
      "10111011000011010011000011111000100111111010011100101101010011011110011000000001111011011101011000101000" when "10000111001",
      "10111011000011010011000011111000100111111010011100101101010011011110011000000001111011011101011000101000" when "10000111010",
      "10111011001001011010001111110101011100010101110011111110100001001001100111010110011100010010001011011100" when "10000111011",
      "10111011001111100001100101001000001111110011110011110111011110010110101110000111110000011000101111010000" when "10000111100",
      "10111011010101101001000011110001011110111001010101100111010100000110000101000111001100100101100010100011" when "10000111101",
      "10111011011011110000101011110001100110001101010101100110100111111111001011100110101011110010001000010000" when "10000111110",
      "10111011100001111000011101001001000010011000110011100011111111000100011111100110011100101101110100100000" when "10000111111",
      "10111011101000000000010111111000010000000110110010110000100010000111010111010001011100110100001101001110" when "10001000000",
      "10111011101000000000010111111000010000000110110010110000100010000111010111010001011100110100001101001110" when "10001000001",
      "10111011101110001000011011111111101100000100011010001100100011011100001001011010110100101101101011011010" when "10001000010",
      "10111011110100010000101001011111110011000000110100110100000110001110110010110000111110110100101000010100" when "10001000011",
      "10111011111010011001000000011001000001101101010001101011100111011000000101111101010100101100110100110100" when "10001000100",
      "10111100000000100001100000101011110100111101000100001100100111110011110100001001110100101001100110111110" when "10001000101",
      "10111100000110101010001010011000101001100101100100010010011000010111111100001000000110001011011001011000" when "10001000110",
      "10111100001100110010111101011111111100011110001110100110100111001101001101110111111001100101001101011000" when "10001000111",
      "10111100001100110010111101011111111100011110001110100110100111001101001101110111111001100101001101011000" when "10001001000",
      "10111100010010111011111010000010001010100000100100101110001110101001010000101101010101000000000101111110" when "10001001001",
      "10111100011001000100111111111111110000101000001101010110000101101010011001111001010111110100000111011000" when "10001001010",
      "10111100011111001110001111011001001011110010110100011111110001110101100001111001110100001101011001001100" when "10001001011",
      "10111100100101010111101000001110111001000000001011101110011010110110000110010111110110001111011001100111" when "10001001100",
      "10111100101011100001001010100001010101010010001010010011011111100000100110111111000111100001101000010100" when "10001001101",
      "10111100101011100001001010100001010101010010001010010011011111100000100110111111000111100001101000010100" when "10001001110",
      "10111100110001101010110110010000111101101100101101011011101100010111101011011001010111000110110010111010" when "10001001111",
      "10111100110111110100101011011110001111010101111000011011110011110100000000011101000101110011000100101110" when "10001010000",
      "10111100111101111110101010001001100111010101110100111101100111101111011011000000010000100110101011100000" when "10001010001",
      "10111101000100001000110010010011100010110110110011001100110100110011001110100010001100100000010010100100" when "10001010010",
      "10111101001010010011000011111100011111000101001010000011111111001010000110000010100001000110101100100100" when "10001010011",
      "10111101010000011101011111000100111001001111010111011001100000110101101101011101001010010010100101100110" when "10001010100",
      "10111101010000011101011111000100111001001111010111011001100000110101101101011101001010010010100101100110" when "10001010101",
      "10111101010110101000000011101101001110100110000000001100101001101000011010000110000100001000101101101000" when "10001010110",
      "10111101011100110010110001110101111100011011110000110010100000100011000000100001011111111001111001000000" when "10001010111",
      "10111101100010111101101001011111100000000101011101000011000110110111000110011000011101000001100100001101" when "10001011000",
      "10111101101001001000101010101010010110111010000000100110011100101101111110101010111101011100111100010001" when "10001011001",
      "10111101101111010011110101010110111110010010011111000001100111010100011111000100101001110100001111000111" when "10001011010",
      "10111101101111010011110101010110111110010010011111000001100111010100011111000100101001110100001111000111" when "10001011011",
      "10111101110101011111001001100101110011101010000100000011111000101011111100111010010111001101011100011001" when "10001011100",
      "10111101111011101010100111010111010100011110000011110011111001000000100000011001111110011100001110100010" when "10001011101",
      "10111110000001110110001110101011111110001101111010111100110001100100111100111000010010111101010011000101" when "10001011110",
      "10111110001000000001111111100100001110011011001110111011011001010100011100101011000110100101000001010110" when "10001011111",
      "10111110001110001101111010000000100010101001101110001011100010111010001111100000000110100001000010000110" when "10001100000",
      "10111110001110001101111010000000100010101001101110001011100010111010001111100000000110100001000010000110" when "10001100001",
      "10111110010100011001111110000001011000011111010000010101001100011111101010000011111110000011100101111000" when "10001100010",
      "10111110011010100110001011100111001101100011110110011001110001000000100101101111001011100101001011001100" when "10001100011",
      "10111110100000110010100010110010011111100001101011000001011011000110101111010000110101011101101101100101" when "10001100100",
      "10111110100110111111000011100011101100000101000010101000011001101011110011010010001101101010110101110001" when "10001100101",
      "10111110101101001011101101111011010000111100011011101100010110000010110111110000010100101011110010010110" when "10001100110",
      "10111110101101001011101101111011010000111100011011101100010110000010110111110000010100101011110010010110" when "10001100111",
      "10111110110011011000100001111001101011111000011110111001101011101001010001001011001110101110000110011101" when "10001101000",
      "10111110111001100101011111011111011010101011111111011001000001011111000010101101100000111000011110001110" when "10001101001",
      "10111110111111110010100110101100111011001011111010111100100101000111011000010000101111010010100000010010" when "10001101010",
      "10111111000101111111110111100010101011001111011010001101100111010001001001100110011000111001100100111111" when "10001101011",
      "10111111001100001101010010000001001000101111110000111001111010000111110101101111010010000100000000011010" when "10001101100",
      "10111111001100001101010010000001001000101111110000111001111010000111110101101111010010000100000000011010" when "10001101101",
      "10111111010010011010110110001000110001101000011110000001010001001101000101101110000011100100101000001001" when "10001101110",
      "10111111011000101000100011111010000011110111001100000011000010111011000110000011111001010001111011000100" when "10001101111",
      "10111111011110110110011011010101011101011011110001001011101011110000000110001001010001000100110011110111" when "10001110000",
      "10111111100101000100011100011011011100011000001111100010010011000011001100110111000001010100100000100101" when "10001110001",
      "10111111101011010010100111001100011110110000110101010110010001100010110001110110110100100110011111000000" when "10001110010",
      "10111111101011010010100111001100011110110000110101010110010001100010110001110110110100100110011111000000" when "10001110011",
      "10111111110001100000111011101001000010101011111101001100111001011100101010110100011111111011011111110110" when "10001110100",
      "10111111110111101111011001110001100110010010001110001111000000010000011100001100100000010101010111000100" when "10001110101",
      "10111111111101111110000001100110100111101110011100010110101010001011111100110110010101000100001111011101" when "10001110110",
      "11000000000100001100110011001000100101001101101000011100110111010010011100001100010100011110010110110100" when "10001110111",
      "11000000000100001100110011001000100101001101101000011100110111010010011100001100010100011110010110110100" when "10001111000",
      "11000000001010011011101110010111111100111111000000100111010010001110011010010101000010111001110001111100" when "10001111001",
      "11000000010000101010110011010101001101010100000000010110000000101110100001110100111100110101111111011000" when "10001111010",
      "11000000010110111010000010000000110100100000010000110001010101101101110010110001101111111001101111101101" when "10001111011",
      "11000000011101001001011010011011010000111001101000110111100101000111001110110011101001000010000111101010" when "10001111100",
      "11000000100011011000111100100101000000111000001101101010111001010101010101110011001001111001000011010110" when "10001111101",
      "11000000100011011000111100100101000000111000001101101010111001010101010101110011001001111001000011010110" when "10001111110",
      "11000000101001101000101000011110100010110110010010011111001010011101100011000101000011000100110010000010" when "10001111111",
      "11000000101111111000011110001000010101010000011001000111110111000111111010111000011101011110000101110001" when "10010000000",
      "11000000110110001000011101100010110110100101010010000101111111000011010111111110001001111001100010000000" when "10010000001",
      "11000000111100011000100110101110100101010101111100110101111111010110101001010010011011101111110110100110" when "10010000010",
      "11000001000010101000111001101100000000000101100111111101110000011110001111100110000001010011110001101111" when "10010000011",
      "11000001000010101000111001101100000000000101100111111101110000011110001111100110000001010011110001101111" when "10010000100",
      "11000001001000111001010110011011100101011001110001011010100101110111101011000100111011000111010001111110" when "10010000101",
      "11000001001111001001111100111101110011111010000110101111001111011010001000111101000010101000101001100000" when "10010000110",
      "11000001010101011010101101010011001010010000100101010001111100011101000001001001000000010111111100111010" when "10010000111",
      "11000001011011101011100111011100000111001001011010011010100000101100010100000110100001100000011000100010" when "10010001000",
      "11000001011011101011100111011100000111001001011010011010100000101100010100000110100001100000011000100010" when "10010001001",
      "11000001100001111100101011011001001001010011000011110000011010101011011001000010001101111110001001010001" when "10010001010",
      "11000001101000001101111001001010101111011110001111011000111100000110001100100101110001001001011101101010" when "10010001011",
      "11000001101110011111010000110001011000011101111100000101010011110001010000010111111001000001111100111011" when "10010001100",
      "11000001110100110000110010001101100011000111011001100000111001011000101011100000100010001010111111101000" when "10010001101",
      "11000001110100110000110010001101100011000111011001100000111001011000101011100000100010001010111111101000" when "10010001110",
      "11000001111011000010011101011111101110010010001000011111011010111110011100100110011001100010010011001111" when "10010001111",
      "11000010000001010100010010101000011000110111111011001011001100001000001101011101110000110101010101110100" when "10010010000",
      "11000010000111100110010001101000000001110100110101010011010110111100111001000011010101111001000111110000" when "10010010001",
      "11000010001101111000011010011111001000000111001100011010001110110010010100000000110010001001111001110111" when "10010010010",
      "11000010010100001010101101001110001010101111101000000011100100101011001000011011001100011110000010010100" when "10010010011",
      "11000010010100001010101101001110001010101111101000000011100100101011001000011011001100011110000010010100" when "10010010100",
      "11000010011010011101001001110101101000110001000010000010111101100101010101001110111101000000001101101110" when "10010010101",
      "11000010100000101111110000010110000001010000100110101010001010011001100001111110111001010010011001010001" when "10010010110",
      "11000010100111000010100000101111110011010101110100110111100001101011010111011111110101001011001111101010" when "10010010111",
      "11000010101101010101011011000011011110001010011110100100011011001011001110001100001100110100101101000010" when "10010011000",
      "11000010101101010101011011000011011110001010011110100100011011001011001110001100001100110100101101000010" when "10010011001",
      "11000010110011101000011111010001100000111010101000110011101101001001100010101110100011101010111100010110" when "10010011010",
      "11000010111001111011101101011010011010110100101100000000001011011100000001110100011100110111111110010001" when "10010011011",
      "11000011000000001111000101011110101011001001010100001011001000010100111011111110001010101001011001100010" when "10010011100",
      "11000011000110100010100111011110110001001011100001001010110111001100110010000010101011100011100100011011" when "10010011101",
      "11000011000110100010100111011110110001001011100001001010110111001100110010000010101011100011100100011011" when "10010011110",
      "11000011001100110110010011011011001100010000100110111001010000111110101011100010000110111111101010001100" when "10010011111",
      "11000011010011001010001001010100011011110000001101100010011010010111100111100011110100110001010000011010" when "10010100000",
      "11000011011001011110001001001010111111000100010001110011001011111000111001100000010111000011110111010011" when "10010100001",
      "11000011011111110010010010111111010101101001000101000111111011101110000010011010001001111001100011111001" when "10010100010",
      "11000011011111110010010010111111010101101001000101000111111011101110000010011010001001111001100011111001" when "10010100011",
      "11000011100110000110100110110001111110111101001101111011001001010110011000001011000111110001111101011110" when "10010100100",
      "11000011101100011011000100100011011010100001100111110100001011000010101011110000000000000011110000000011" when "10010100101",
      "11000011110010101111101100010100000111111001100011110101111101000110111111011101011001011011100100011011" when "10010100110",
      "11000011111001000100011110000100100110101010101000101101110011000000111110101101011001000000111011111000" when "10010100111",
      "11000011111001000100011110000100100110101010101000101101110011000000111110101101011001000000111011111000" when "10010101000",
      "11000011111111011001011001110101010110011100110011000010001010010011001000010111100101010101100010000010" when "10010101001",
      "11000100000101101110011111100110110110111010010101100001011111010100111101001000011011111100011011101001" when "10010101010",
      "11000100001100000011101111011001100111101111111001010001000011111000100011001111110000010110000100100110" when "10010101011",
      "11000100010010011001001001001110001000101100011101111011110111100101110001000001001011100010111011111001" when "10010101100",
      "11000100010010011001001001001110001000101100011101111011110111100101110001000001001011100010111011111001" when "10010101101",
      "11000100011000101110101101000100111001100001011010000001100010001011001111100100100100101010010000100010" when "10010101110",
      "11000100011111000100011010111110011010000010011011000101001111100101100111010111001100110011101001001000" when "10010101111",
      "11000100100101011010010010111011001010000101100101111100101101111101001000000001101010111010011110111110" when "10010110000",
      "11000100101011110000010100111011101001100011010110111111001101011001111101001001100111000000101000000110" when "10010110001",
      "11000100101011110000010100111011101001100011010110111111001101011001111101001001100111000000101000000110" when "10010110010",
      "11000100110010000110100001000000011000010110100010010100100001101111100001101001001000001010111000100001" when "10010110011",
      "11000100111000011100110111001001110110011100010100000100000101111111000011011001001100011110000011100011" when "10010110100",
      "11000100111110110011010111011000100011110100010000100100000001110001101000111111000111000110000010101101" when "10010110101",
      "11000101000101001010000001101101000000100000010100101000010000101010001011010000010110001010101010000001" when "10010110110",
      "11000101000101001010000001101101000000100000010100101000010000101010001011010000010110001010101010000001" when "10010110111",
      "11000101001011100000110110000111101100100100110101110001101011001111010100100011000111110111000000000001" when "10010111000",
      "11000101010001110111110100101001001000001000100010011101010010001101110111100101001101000000110110010110" when "10010111001",
      "11000101011000001110111101010001110011010100100010010011011011010011101111110101011110101101100100011000" when "10010111010",
      "11000101011110100110010000000010001110010100010110010111000000000011111101100000000100001001110010100000" when "10010111011",
      "11000101011110100110010000000010001110010100010110010111000000000011111101100000000100001001110010100000" when "10010111100",
      "11000101100100111101101100111010111001010101111001010100101110100011101110111111101110101000100010101100" when "10010111101",
      "11000101101011010101010011111100010100101001011111110010011100000001001010001010101010100101111010110010" when "10010111110",
      "11000101110001101101000101000111000000100001111000011110011001010011100111010011101110011000101111011000" when "10010111111",
      "11000101110001101101000101000111000000100001111000011110011001010011100111010011101110011000101111011000" when "10011000000",
      "11000101111000000101000000011011011101010100001100011110101001010110010000001100011001110110010100100110" when "10011000001",
      "11000101111110011101000101111010001011010111111111100000011001011100110101010111000100101011010101010000" when "10011000010",
      "11000110000100110101010101100011101011000111010000000111011011100011001011111100000101010101001001001011" when "10011000011",
      "11000110001011001101101111011000011100111110010111111101100010010111100110010111100110011000000011110100" when "10011000100",
      "11000110001011001101101111011000011100111110010111111101100010010111100110010111100110011000000011110100" when "10011000101",
      "11000110010001100110010011011001000001011100001100000001111111100000011010011001001101001000100011100100" when "10011000110",
      "11000110010111111111000001100101111001000001111100111001000011011101000110110001100010000000010011000010" when "10011000111",
      "11000110011110010111111001111111100100010011010110111011011111100011001011001101011001000011011000101100" when "10011001000",
      "11000110100100110000111100100110100011110110100010100110001001110111000101000001001000001111000111111100" when "10011001001",
      "11000110100100110000111100100110100011110110100010100110001001110111000101000001001000001111000111111100" when "10011001010",
      "11000110101011001010001001011011011000010100000100101001100011000001100011001010001000001001110010000111" when "10011001011",
      "11000110110001100011100000011110100010010110111110011001011110000001100100001111101100010010011111010100" when "10011001100",
      "11000110110111111101000001110000100010101100101101111100101001111011010001001111110000100001101000000000" when "10011001101",
      "11000110110111111101000001110000100010101100101101111100101001111011010001001111110000100001101000000000" when "10011001110",
      "11000110111110010110101101010001111010000101001110011100011101100100000111100111001011000101001001111110" when "10011001111",
      "11000111000100110000100011000011001001010010111000010100100101001100100101101000100100001001001111000000" when "10011010000",
      "11000111001011001010100011000100110001001010100001100010110010000111101011111000000111001100011011100000" when "10011010001",
      "11000111010001100100101101010111010010100011011101110110101100010000100110100101110101011000000111000111" when "10011010010",
      "11000111010001100100101101010111010010100011011101110110101100010000100110100101110101011000000111000111" when "10011010011",
      "11000111010111111111000001111011001110010111011111000001100101101110110010000011010100011001000101100001" when "10011010100",
      "11000111011110011001100000110001000101100010110101000110010000011000101100110101001010000010101000001010" when "10011010101",
      "11000111100100110100001001111001011001000100001110101000110101010101101011000011101001111110101111000101" when "10011010110",
      "11000111100100110100001001111001011001000100001110101000110101010101101011000011101001111110101111000101" when "10011010111",
      "11000111101011001110111101010100101001111100111000111110101110011110111101110001110001010001111111011011" when "10011011000",
      "11000111110001101001111011000011011001010000100000011110100010000000100001100100100010000111110011110000" when "10011011001",
      "11000111111000000101000011000110001000000101010000101111111111111001100111101000101001010101011110001110" when "10011011010",
      "11000111111110100000010101011101010111100011110100111100000001011101101100100111001111100111001001101010" when "10011011011",
      "11000111111110100000010101011101010111100011110100111100000001011101101100100111001111100111001001101010" when "10011011100",
      "11001000000100111011110010001001101000110111010111111100101010110101110000011110010000111010010101011000" when "10011011101",
      "11001000001011010111011001001011011101001101100100101101001110100010100010110100001110000100111010011110" when "10011011110",
      "11001000010001110011001010100011010101110110100110011010010010111111110111000010100110101111101010011000" when "10011011111",
      "11001000010001110011001010100011010101110110100110011010010010111111110111000010100110101111101010011000" when "10011100000",
      "11001000011000001111000110010001110100000101001000110001111010001001010011110101100100011110001110111100" when "10011100001",
      "11001000011110101011001100010111011001001110011000010011101011000000110001100010111011011110001111000011" when "10011100010",
      "11001000100101000111011100110100100110101010000010100000111101010110111010111110000001100010100000101000" when "10011100011",
      "11001000100101000111011100110100100110101010000010100000111101010110111010111110000001100010100000101000" when "10011100100",
      "11001000101011100011110111101001111101110010010110001101000111010110000100010001011000100111101101000010" when "10011100101",
      "11001000110010000000011100111000000000000100000011101101101101001111101011101010101000000011101000000101" when "10011100110",
      "11001000111000011101001100011111001110111110011101001010110011001100110111101000011101110001111111110100" when "10011100111",
      "11001000111110111010000110100000001100000011010110101111010001000010000110011110001111101111000100101000" when "10011101000",
      "11001000111110111010000110100000001100000011010110101111010001000010000110011110001111101111000100101000" when "10011101001",
      "11001001000101010111001010111011011000110111000110111001001000000110100011000011110101011011100000010100" when "10011101010",
      "11001001001011110100011001110001010111000000100110101001111011001111010010101100010001111100110011101011" when "10011101011",
      "11001001010010010001110011000010101000001001010001110111001000101110110000000001000111110011000011110011" when "10011101100",
      "11001001010010010001110011000010101000001001010001110111001000101110110000000001000111110011000011110011" when "10011101101",
      "11001001011000101111010110101111101101111101000111011010100110011000100111000011110001101111010000100000" when "10011101110",
      "11001001011111001101000100111001001010001010101001100010111111101010100110011001111110010110000011011110" when "10011101111",
      "11001001100101101010111101011111011110100010111110000100010101111010011001101101101111001000110000101000" when "10011110000",
      "11001001100101101010111101011111011110100010111110000100010101111010011001101101101111001000110000101000" when "10011110001",
      "11001001101100001001000000100011001100111001101110101000100010101001000001101101000000001010100011101000" when "10011110010",
      "11001001110010100111001110000100110111000101001000111111111011111011111101111000100001100010000010011000" when "10011110011",
      "11001001111001000101100110000100111110111101111111010001111010111100011100010101010001101111100111000011" when "10011110100",
      "11001001111111100100001000100100000110011111101000001101100100011101000011110111001101111000001100000110" when "10011110101",
      "11001001111111100100001000100100000110011111101000001101100100011101000011110111001101111000001100000110" when "10011110110",
      "11001010000110000010110101100010101111100111111111011010010011100110001100111111110011011001000001100110" when "10011110111",
      "11001010001100100001101101000001011100010111100101101000100110101001011110001110010110111101110001100001" when "10011111000",
      "11001010010011000000101111000000101110110001100001000010101101111100100000000011111100000101000001101100" when "10011111001",
      "11001010010011000000101111000000101110110001100001000010101101111100100000000011111100000101000001101100" when "10011111010",
      "11001010011001011111111011100001001000111011011101011101011100111011011101100000000010000001110001100010" when "10011111011",
      "11001010011111111111010010100011001100111101101100101000111101010011100101011111000100111001110010001000" when "10011111100",
      "11001010100110011110110100000111011101000011000110100001100100010110000010000111011011100001110010011001" when "10011111101",
      "11001010100110011110110100000111011101000011000110100001100100010110000010000111011011100001110010011001" when "10011111110",
      "11001010101100111110100000001110011011011001001001100000101010010011011010010101000110101000111011111011" when "10011111111",
      "11001010110011011110010110111000101010001111111010101101100100000000010010111000010001100101001111111010" when "10100000000",
      "11001010111001111110011000000110101011111010000110001110011110100011000011011110010001100011000011101000" when "10100000001",
      "11001010111001111110011000000110101011111010000110001110011110100011000011011110010001100011000011101000" when "10100000010",
      "11001011000000011110100011111001000010101100111111011001011101001011010101000000011101111001110010101010" when "10100000011",
      "11001011000110111110111010010000010001000000100001000101011001010011011101111000001010011001000101110110" when "10100000100",
      "11001011001101011111011011001100111001001111001101111011000100101100010001011010011011000010010100010100" when "10100000101",
      "11001011001101011111011011001100111001001111001101111011000100101100010001011010011011000010010100010100" when "10100000110",
      "11001011010100000000000110101111011101110110010000100110001101110011010111100010011001010100010010011100" when "10100000111",
      "11001011011010100000111100111000100001010101011100000110100110010100100001110100100010110001100100011111" when "10100001000",
      "11001011100001000001111101101000100110001111001100000001001011110110010011001000111010011101001011000011" when "10100001001",
      "11001011100001000001111101101000100110001111001100000001001011110110010011001000111010011101001011000011" when "10100001010",
      "11001011100111100011001001000000001111001000100100110001010010110010001111001110011000101110001010001010" when "10100001011",
      "11001011101110000100011110111111111110101001010011111001110011011001000111011100100111110000101011001101" when "10100001100",
      "11001011110100100101111111101000010111011011110000010110011001000011011010001110001110110010011001101111" when "10100001101",
      "11001011110100100101111111101000010111011011110000010110011001000011011010001110001110110010011001101111" when "10100001110",
      "11001011111011000111101010111001111100001100111010101100110011101110011010100000100010010001100110111111" when "10100001111",
      "11001100000001101001100000110101001111101100011101011110001011100110010100111010000100110001000010111100" when "10100010000",
      "11001100001000001011100001011010110100101100101101011000010110111101100111111100111001101111111111001110" when "10100010001",
      "11001100001000001011100001011010110100101100101101011000010110111101100111111100111001101111111111001110" when "10100010010",
      "11001100001110101101101100101011001110000010101001100111010010010010000101001101100010110101000011101100" when "10100010011",
      "11001100010101010000000010100110111110100101111100000110011010011111110000111011010110111100001010000101" when "10100010100",
      "11001100011011110010100011001110101001010000111001110010001001100010010101111010111011101100001000110111" when "10100010101",
      "11001100011011110010100011001110101001010000111001110010001001100010010101111010111011101100001000110111" when "10100010110",
      "11001100100010010101001110100010110001000000100010111001010101000101000011100111000001111111111000010000" when "10100010111",
      "11001100101000111000000100100011111000110100100011001110101111100001101100000000100001001000011101011001" when "10100011000",
      "11001100101111011011000101010010100011101111010010011010101011001110110111101001100101111011001111010010" when "10100011001",
      "11001100101111011011000101010010100011101111010010011010101011001110110111101001100101111011001111010010" when "10100011010",
      "11001100110101111110010000101111010100110101110100001100011111111110000101011100100111011111000101111000" when "10100011011",
      "11001100111100100001100110111010101111001111111000101100010010101001101100100010101111000000000000000110" when "10100011100",
      "11001101000011000101000111110101010110000111111100101100011111010011010110010010011101010111110101010100" when "10100011101",
      "11001101000011000101000111110101010110000111111100101100011111010011010110010010011101010111110101010100" when "10100011110",
      "11001101001001101000110011011111101100101011001001111011100101010011000110100010010111010110100111010000" when "10100011111",
      "11001101010000001100101001111010010110001001010111010101110101110111101000011111111111100100001011110100" when "10100100000",
      "11001101010110110000101011000101110101110101001001010111000100110111110110011111000101011000111010001111" when "10100100001",
      "11001101010110110000101011000101110101110101001001010111000100110111110110011111000101011000111010001111" when "10100100010",
      "11001101011101010100110111000010101111000011110010001100011011110110010010111001010000000011010101010001" when "10100100011",
      "11001101100011111001001101110001100101001101010010000110001111010110101000111010001110011101100010101101" when "10100100100",
      "11001101101010011101101111010010111011101100010111101001110110100101101011011000110110010110101011010100" when "10100100101",
      "11001101101010011101101111010010111011101100010111101001110110100101101011011000110110010110101011010100" when "10100100110",
      "11001101110001000010011011100111010101111110100000000011100101010100001000100001000000001011101000111010" when "10100100111",
      "11001101110111100111010010101111010111100011110111011000101000000100101000110110110000110101111111010100" when "10100101000",
      "11001101111110001100010100101011100011111111011000111001000010101101010000011111000110111001001101000011" when "10100101001",
      "11001101111110001100010100101011100011111111011000111001000010101101010000011111000110111001001101000011" when "10100101010",
      "11001110000100110001100001011100011110110110101111010001110001001100111000111110100110001101010101100011" when "10100101011",
      "11001110001011010110111001000010101011110010010100111110101010110100111011000010100011010010101100111100" when "10100101100",
      "11001110010001111100011011011110101110011101010100011100100111100111011110101101010110011100110010001100" when "10100101101",
      "11001110010001111100011011011110101110011101010100011100100111100111011110101101010110011100110010001100" when "10100101110",
      "11001110011000100010001000110001001010100101101000011011101000001010101001000010100110111011010011000000" when "10100101111",
      "11001110011111001000000000111010100011111011111100010000111111110000111110010100000110110111011010101100" when "10100110000",
      "11001110011111001000000000111010100011111011111100010000111111110000111110010100000110110111011010101100" when "10100110001",
      "11001110100101101110000011111011011110010011101100001001100000110111101111110100100010100000110110110100" when "10100110010",
      "11001110101100010100010001110100011101100011000101011011101011111011001100011001001111100010110110000100" when "10100110011",
      "11001110110010111010101010100110000101100011000110111010000000100001001010111000010100101100011100000101" when "10100110100",
      "11001110110010111010101010100110000101100011000110111010000000100001001010111000010100101100011100000101" when "10100110101",
      "11001110111001100001001110010000111010001111100001000101010000111010100101110100101110000010000110000010" when "10100110110",
      "11001111000000000111111100110101011111100110110110011110110111111011111111101101111111010000010001101101" when "10100110111",
      "11001111000110101110110110010100011001101010011011111011010001001101100111001101110011010000010011101101" when "10100111000",
      "11001111000110101110110110010100011001101010011011111011010001001101100111001101110011010000010011101101" when "10100111001",
      "11001111001101010101111010101110001100011110011000110100010011110011010010110001010111000001110011110000" when "10100111010",
      "11001111010011111101001010000011011100001001100111011011101111001100101011010001001101100100001101011110" when "10100111011",
      "11001111011010100100100100010100101100110101110101001101101010101101111101001110001010111101000110100111" when "10100111100",
      "11001111011010100100100100010100101100110101110101001101101010101101111101001110001010111101000110100111" when "10100111101",
      "11001111100001001100001001100010100010101111100011000011000111010001101000001110010110010001110100010101" when "10100111110",
      "11001111100111110011111001101101100010000110000101100100100011100011100100011001100100001100110111100110" when "10100111111",
      "11001111100111110011111001101101100010000110000101100100100011100011100100011001100100001100110111100110" when "10101000000",
      "11001111101110011011110100110110001111001011100101011100100010100101110101101000101111010010110111101111" when "10101000001",
      "11001111110101000011111010111101001110010100111111101010010100101111100100100000000111001110100000010110" when "10101000010",
      "11001111111011101100001100000011000011111010000101110100100011000110010100110000100100111000010010100100" when "10101000011",
      "11001111111011101100001100000011000011111010000101110100100011000110010100110000100100111000010010100100" when "10101000100",
      "11010000000010010100101000001000010100010101011110011011111101010010010001100000100111010101011101001110" when "10101000101",
      "11010000001000111101001111001101100100000100100101001110001001101101100111000001110100011001011001110110" when "10101000110",
      "11010000001111100110000001010011010111100111101011011000011000001111100010011100001110111111001100001110" when "10101000111",
      "11010000001111100110000001010011010111100111101011011000011000001111100010011100001110111111001100001110" when "10101001000",
      "11010000010110001110111110011010010011100001110111111010010111010011001111011101001110010100100001111111" when "10101001001",
      "11010000011100111000000110100010111100011001000111111001001011011011001100011011111010001110000000101110" when "10101001010",
      "11010000011100111000000110100010111100011001000111111001001011011011001100011011111010001110000000101110" when "10101001011",
      "11010000100011100001011001101101110110110110001110110010001001010001001101001001101011010100111101011000" when "10101001100",
      "11010000101010001010110111111011100111100100110110101101110010000011100100101001101001010010101111110100" when "10101001101",
      "11010000110000110100100001001100110011010011100000110010110010011111101110101110011101001011100101010010" when "10101001110",
      "11010000110000110100100001001100110011010011100000110010110010011111101110101110011101001011100101010010" when "10101001111",
      "11010000110111011110010101100001111110110011100101011001000100001010110001100010001011100100001010011110" when "10101010000",
      "11010000111110001000010100111011101110111001010100011100110001011000010000000000100111110010001111111101" when "10101010001",
      "11010000111110001000010100111011101110111001010100011100110001011000010000000000100111110010001111111101" when "10101010010",
      "11010001000100110010011111011010101000011011110101110001011011011111100101110000110000111000010111011010" when "10101010011",
      "11010001001011011100110100111111010000010101001001010101000011110000100101001110101000101000110011111100" when "10101010100",
      "11010001010010000111010101101010001011100010000111100011010110100111010000111011010110000100000000101000" when "10101010101",
      "11010001010010000111010101101010001011100010000111100011010110100111010000111011010110000100000000101000" when "10101010110",
      "11010001011000110010000001011011111111000010100001101000111001011111101000101101100110011010010101110110" when "10101010111",
      "11010001011111011100111000010101001111111001000001110110011011001001100100000001100010101010000100110100" when "10101011000",
      "11010001100110000111111010010110100011001011001011110100000110011101010010001011010010111111000111110011" when "10101011001",
      "11010001100110000111111010010110100011001011001011110100000110011101010010001011010010111111000111110011" when "10101011010",
      "11010001101100110011000111100000011110000001011100110100110111110000111001110100001110100100010011001001" when "10101011011",
      "11010001110011011110011111110011100101100111001100001001110100101111010000101111011011011100110100101111" when "10101011100",
      "11010001110011011110011111110011100101100111001100001001110100101111010000101111011011011100110100101111" when "10101011101",
      "11010001111010001010000011010000011111001010101011010101100110110000100101010110101001000001000101000001" when "10101011110",
      "11010010000000110101110001110111101111111101000110011111110111110101010011000101010110111011100010100000" when "10101011111",
      "11010010000111100001101011101001111101010010100100101000110010000011011011001100100011000010010111001100" when "10101100000",
      "11010010000111100001101011101001111101010010100100101000110010000011011011001100100011000010010111001100" when "10101100001",
      "11010010001110001101110000100111101100100010000111111100100001100110111011011110000010000111101011010010" when "10101100010",
      "11010010010100111010000000110001100011000101101110000110111001010101011100010011010001110110011010001100" when "10101100011",
      "11010010010100111010000000110001100011000101101110000110111001010101011100010011010001110110011010001100" when "10101100100",
      "11010010011011100110011100001000000110011010010000100110111001110101101111110111111101101011101011100111" when "10101100101",
      "11010010100010010011000010101011111011111111100101000010011011001011011100000101011100110101101001100001" when "10101100110",
      "11010010101000111111110100011101101001011000011101011001111001000111001001000000111100111000011011110011" when "10101100111",
      "11010010101000111111110100011101101001011000011101011001111001000111001001000000111100111000011011110011" when "10101101000",
      "11010010101111101100110001011101110100001010101000011100000001111011101101110010111010110000101010100000" when "10101101001",
      "11010010110110011001111001101101000001111110110001111001100111111000110101110010111011100001010101111110" when "10101101010",
      "11010010110110011001111001101101000001111110110001111001100111111000110101110010111011100001010101111110" when "10101101011",
      "11010010111101000111001101001011111000100000100010111001010101001011011000001000000110010000101000100011" when "10101101100",
      "11010011000011110100101011111010111101011110100010001011100010100011111011100010110010001100101110000100" when "10101101101",
      "11010011001010100010010101111010110110101010010100011110010000100100000000111001001110000111101010100011" when "10101101110",
      "11010011001010100010010101111010110110101010010100011110010000100100000000111001001110000111101010100011" when "10101101111",
      "11010011010001010000001011001100001001111000011100110001000011010010001110010101011001101111001000000011" when "10101110000",
      "11010011010111111110001011101111011101000000011100101001000000110101110101100111011101111011010101110100" when "10101110001",
      "11010011010111111110001011101111011101000000011100101001000000110101110101100111011101111011010101110100" when "10101110010",
      "11010011011110101100010111100101010101111100110100100100110010011010001111110100100110001000000101000001" when "10101110011",
      "11010011100101011010101110101110011010101011000100010000100111111010101000111111010011100010100010110010" when "10101110100",
      "11010011100101011010101110101110011010101011000100010000100111111010101000111111010011100010100010110010" when "10101110101",
      "11010011101100001001010001001011010001001011101010111010011110010110010110001010111010010000110010011001" when "10101110110",
      "11010011110010110111111110111100011111100010000111100110001000101110010000100000110000110010001101010010" when "10101110111",
      "11010011111001100110111000000010101011110100111001100001011011101011110000000010110011110101011111011000" when "10101111000",
      "11010011111001100110111000000010101011110100111001100001011011101011110000000010110011110101011111011000" when "10101111001",
      "11010100000000010101111100011110011100001101100000011000011011110001100000111011111010111111000110111110" when "10101111010",
      "11010100000111000101001100010000010110111000011100101001101110010110101110000011010101111100011100101001" when "10101111011",
      "11010100000111000101001100010000010110111000011100101001101110010110101110000011010101111100011100101001" when "10101111100",
      "11010100001101110100100111011001000010000101001111111010101101001100111011101101100111000011000100000110" when "10101111101",
      "11010100010100100100001101111001000100000110011101001011111100110001001101101010001101000001101111100010" when "10101111110",
      "11010100011011010011111111110001000011010001101001001101100101001000110011010010001100110010000110001101" when "10101111111",
      "11010100011011010011111111110001000011010001101001001101100101001000110011010010001100110010000110001101" when "10110000000",
      "11010100100010000011111101000001100101111111011010110011101101101001110101010001001011100101110010101110" when "10110000001",
      "11010100101000110100000101101011010010101011011011001010111011010000011111110110101010111010001110011001" when "10110000010",
      "11010100101000110100000101101011010010101011011011001010111011010000011111110110101010111010001110011001" when "10110000011",
      "11010100101111100100011001101110101111110100010110001100110001100001000101000011011000110000111101110000" when "10110000100",
      "11010100110110010100111001001100100011111011111010110100010110010111010010001010101010100010101101011111" when "10110000101",
      "11010100110110010100111001001100100011111011111010110100010110010111010010001010101010100010101101011111" when "10110000110",
      "11010100111101000101100100000101010101100110111011010010111000100011010100000101011011111110001000100110" when "10110000111",
      "11010101000011110110011010011001101011011101001101100100011000110101000101111001010001000100000110110110" when "10110001000",
      "11010101001010100111011100001010001100001001101011100100010101110110000101011010111111110111100111101010" when "10110001001",
      "11010101001010100111011100001010001100001001101011100100010101110110000101011010111111110111100111101010" when "10110001010",
      "11010101010001011000101001010111011110011010010011100010011010110010001001011001101110000001100000100001" when "10110001011",
      "11010101011000001010000010000010001001000000001000010111010000101111110101000011110110010111000111100010" when "10110001100",
      "11010101011000001010000010000010001001000000001000010111010000101111110101000011110110010111000111100010" when "10110001101",
      "11010101011110111011100110001010110010101111010001111001010010111000100100111101010100000111100011111011" when "10110001110",
      "11010101100101101101010101110010000010011110111101010001100101010001010001000010111011101101011111000110" when "10110001111",
      "11010101100101101101010101110010000010011110111101010001100101010001010001000010111011101101011111000110" when "10110010000",
      "11010101101100011111010000111000011111001001011101010000101110100011011111111100010100100011100001101010" when "10110010001",
      "11010101110011010001010111011110101111101100001010100011110100011000000111100010110100000000001010011001" when "10110010010",
      "11010101111010000011101001100101011011000111100100001001011010100011010111001001000111001010110001010000" when "10110010011",
      "11010101111010000011101001100101011011000111100100001001011010100011010111001001000111001010110001010000" when "10110010100",
      "11010110000000110110000111001101001000011111001111100110100101000011000111010100101000001111011110110010" when "10110010101",
      "11010110000111101000110000010110011110111001111001011011111100101111101011111110101011110010011011011100" when "10110010110",
      "11010110000111101000110000010110011110111001111001011011111100101111101011111110101011110010011011011100" when "10110010111",
      "11010110001110011011100101000010000101100001010101011010110110111111100100111001000011100101001000101100" when "10110011000",
      "11010110010101001110100101010000100011100010011110111010011111111110101001010110100110101010101010010100" when "10110011001",
      "11010110010101001110100101010000100011100010011110111010011111111110101001010110100110101010101010010100" when "10110011010",
      "11010110011100000001110001000010100000001101011001001101000111111001001011011110000001101000110010001100" when "10110011011",
      "11010110100010110101001000011000100010110101001111110101010010111011001111110010000110011110010011000101" when "10110011100",
      "11010110100010110101001000011000100010110101001111110101010010111011001111110010000110011110010011000101" when "10110011101",
      "11010110101001101000101011010011010010110000010110111011001100000100110110000000001000111000101100001101" when "10110011110",
      "11010110110000011100011001110011010111011000001011100001111010110011001111101010101010101110010101010100" when "10110011111",
      "11010110110111010000010011111001011000001001010011111100111011100000000001101011110011110110000110100011" when "10110100000",
      "11010110110111010000010011111001011000001001010011111100111011100000000001101011110011110110000110100011" when "10110100001",
      "11010110111110000100011001100101111100100011100000000101011010110110001101110000001001110010010110100111" when "10110100010",
      "11010111000100111000101010111001101100001001101001101111110011111110000000110000010101101011101001011000" when "10110100011",
      "11010111000100111000101010111001101100001001101001101111110011111110000000110000010101101011101001011000" when "10110100100",
      "11010111001011101101000111110101001110100001110101000001010001011111100011010101000010000111111000000110" when "10110100101",
      "11010111010010100001110000011001001011010101010000100101010001011101001001110110010111000100101110010011" when "10110100110",
      "11010111010010100001110000011001001011010101010000100101010001011101001001110110010111000100101110010011" when "10110100111",
      "11010111011001010110100100100110001010010000010110000011001100000101100001001101010111100000111100000100" when "10110101000",
      "11010111100000001011100100011100110011000010101010010011111101011110010101110011100011001111001001110110" when "10110101001",
      "11010111100000001011100100011100110011000010101010010011111101011110010101110011100011001111001001110110" when "10110101010",
      "11010111100111000000101111111101101101011110111101110111110010000111110010010001111111000110111101001001" when "10110101011",
      "11010111101101110110000111001001100001011011001101001011110110011001010011100111000111001110001010011101" when "10110101100",
      "11010111101101110110000111001001100001011011001101001011110110011001010011100111000111001110001010011101" when "10110101101",
      "11010111110100101011101010000000110110110000100001000000001000111000010000001111110000100100111001001100" when "10110101110",
      "11010111111011100001011000100100010101011011001110101101001111101000110000000101100011011011010101100110" when "10110101111",
      "11010111111011100001011000100100010101011011001110101101001111101000110000000101100011011011010101100110" when "10110110000",
      "11011000000010010111010010110100100101011010111000101010010000011001010011001010011100000000100010100101" when "10110110001",
      "11011000001001001101011000110010001110110010001110100010101011101001100100111110100101001110000111001010" when "10110110010",
      "11011000010000000011101010011101111001100111001101101100011010101100111010100011100111110110000001000000" when "10110110011",
      "11011000010000000011101010011101111001100111001101101100011010101100111010100011100111110110000001000000" when "10110110100",
      "11011000010110111010000111111000001110000011000001011101110000101000111001010101110001000101101010100111" when "10110110101",
      "11011000011101110000110001000001110100010010000011100011011110010000100101001000111100101100110010100111" when "10110110110",
      "11011000011101110000110001000001110100010010000011100011011110010000100101001000111100101100110010100111" when "10110110111",
      "11011000100100100111100101111011010100100011111100010110111000111100110011011101111001011111001101001000" when "10110111000",
      "11011000101011011110100110100101010111001011100011010100000100100010000010101000101010111111000010011001" when "10110111001",
      "11011000101011011110100110100101010111001011100011010100000100100010000010101000101010111111000010011001" when "10110111010",
      "11011000110010010101110011000000100100011110111111010000000000000100010011000111111000000001011001100000" when "10110111011",
      "11011000111001001101001011001101100100110111100110101110110101101001100001110001100100010010001111100101" when "10110111100",
      "11011000111001001101001011001101100100110111100110101110110101101001100001110001100100010010001111100101" when "10110111101",
      "11011001000000000100101111001101000000110010000000011010001101001011000001100000100010011101100011000110" when "10110111110",
      "11011001000110111100011110111111100000101110000011010111100010000110010011010010011101010100001110011110" when "10110111111",
      "11011001000110111100011110111111100000101110000011010111100010000110010011010010011101010100001110011110" when "10111000000",
      "11011001001101110100011010100101101101001110110111011110011100001101111011001101001000000010101100110000" when "10111000001",
      "11011001010100101100100010000000001110111010110101101111001011011010110001100110111001011110000100110011" when "10111000010",
      "11011001010100101100100010000000001110111010110101101111001011011010110001100110111001011110000100110011" when "10111000011",
      "11011001011011100100110101001111101110011011101000101001000110011110001111010100001010001011101011111110" when "10111000100",
      "11011001100010011101010100010100110100011110001100100001001100110101110100000001100011010101101101110001" when "10111000101",
      "11011001100010011101010100010100110100011110001100100001001100110101110100000001100011010101101101110001" when "10111000110",
      "11011001101001010101111111010000001001110010101111111000101011100000100110001000100010111110111100110001" when "10111000111",
      "11011001110000001110110110000010010111001100110011110011100100110111001011010001110010110111110110100100" when "10111001000",
      "11011001110000001110110110000010010111001100110011110011100100110111001011010001110010110111110110100100" when "10111001001",
      "11011001110111000111111000101100000101100011001100001111011011100110011000111110101000011000001010100010" when "10111001010",
      "11011001111110000001000111001101111101110000000000011010000000101101011100111000111110110010110000010010" when "10111001011",
      "11011001111110000001000111001101111101110000000000011010000000101101011100111000111110110010110000010010" when "10111001100",
      "11011010000100111010100001101000101000110000101011001000000100011111111100001110111001011101011111000011" when "10111001101",
      "11011010001011110100000111111100101111100101111011001100001010101100001010000100111000011100111001110001" when "10111001110",
      "11011010001011110100000111111100101111100101111011001100001010101100001010000100111000011100111001110001" when "10111001111",
      "11011010010010101101111010001010111011010011110011101101100001100110010100010000001001001011110110010110" when "10111010000",
      "11011010011001100111111000010011110101000001101100011110111100011001000110101111111100010001111110000001" when "10111010001",
      "11011010011001100111111000010011110101000001101100011110111100011001000110101111111100010001111110000001" when "10111010010",
      "11011010100000100010000010011000000101111010010010010101110000011100000101100011001011001001110101000101" when "10111010011",
      "11011010100111011100011000011000010111001011100111100000110101110000011100111101011010011000010101101001" when "10111010100",
      "11011010101110010110111010010101010010000111000011111111101010100100101000100100101001101011100111000111" when "10111010101",
      "11011010101110010110111010010101010010000111000011111111101010100100101000100100101001101011100111000111" when "10111010110",
      "11011010110101010001101000001111100000000001010101111001011001111111010001000111000111011111110000010010" when "10111010111",
      "11011010111100001100100010000111101010010010100001110100000101110010000001011110100100100100011111011110" when "10111011000",
      "11011010111100001100100010000111101010010010100001110100000101110010000001011110100100100100011111011110" when "10111011001",
      "11011011000011000111100111111110011010010110000011001011110011010100110011011100101011101111100000000010" when "10111011010",
      "11011011001010000010111001110100011001101010101100101001111011101001110100100010001011001101000011110010" when "10111011011",
      "11011011001010000010111001110100011001101010101100101001111011101001110100100010001011001101000011110010" when "10111011100",
      "11011011010000111110010111101010010001110010101000011100011110101011000011101000100110111011011101000110" when "10111011101",
      "11011011010111111010000001100000101100010011011000101101011001100001101000001100110111101101111001011011" when "10111011110",
      "11011011010111111010000001100000101100010011011000101101011001100001101000001100110111101101111001011011" when "10111011111",
      "11011011011110110101110111011000010010110101110111111010000000000111100011101110100111011001101111110010" when "10111100000",
      "11011011100101110001111001010001101111000110011001001010011001110100011110011111001001001101000001000010" when "10111100001",
      "11011011100101110001111001010001101111000110011001001010011001110100011110011111001001001101000001000010" when "10111100010",
      "11011011101100101110000111001101101010110100101000101001000001010101110000100000011100111111101100001100" when "10111100011",
      "11011011101100101110000111001101101010110100101000101001000001010101110000100000011100111111101100001100" when "10111100100",
      "11011011110011101010100001001100101111110011101011111010000111110010100111111011011101011010101111010001" when "10111100101",
      "11011011111010100111000111001111100111111010000010010011011010111100101101111010101011010000000110100110" when "10111100110",
      "11011011111010100111000111001111100111111010000010010011011010111100101101111010101011010000000110100110" when "10111100111",
      "11011100000001100011111001010110111101000001100101010011101110101101101011011100111100010110110010100100" when "10111101000",
      "11011100001000100000110111100011011001000111101000111010101001110010001111011010001001101101110000101010" when "10111101001",
      "11011100001000100000110111100011011001000111101000111010101001110010001111011010001001101101110000101010" when "10111101010",
      "11011100001111011110000001110101100110001100111100000000010101100011010111011010001110101111111111010000" when "10111101011",
      "11011100010110011011011000001110001110010101101000101101010001001101111101000101000100000100001001011011" when "10111101100",
      "11011100010110011011011000001110001110010101101000101101010001001101111101000101000100000100001001011011" when "10111101101",
      "11011100011101011000111010101101111011101001010100110010001000001001101001011000011001001011001110001001" when "10111101110",
      "11011100100100010110101001010101011000010011000001111111101011011111001111110111001011100011010011001010" when "10111101111",
      "11011100100100010110101001010101011000010011000001111111101011011111001111110111001011100011010011001010" when "10111110000",
      "11011100101011010100100100000101001110100001001110011110101110111111010011101100010101011111001100011101" when "10111110001",
      "11011100110010010010101010111110001000100101110101001000001001001001011000100001001100111000101100010101" when "10111110010",
      "11011100110010010010101010111110001000100101110101001000001001001001011000100001001100111000101100010101" when "10111110011",
      "11011100111001010000111110000000110000110110001101111100110110100100100001001110101001000010100011010000" when "10111110100",
      "11011101000000001111011101001101110001101011001110011110000000101001011110110110000110111001000111111100" when "10111110101",
      "11011101000000001111011101001101110001101011001110011110000000101001011110110110000110111001000111111100" when "10111110110",
      "11011101000111001110001000100101110101100001001010000101000111011111010001110110100101000101000101110111" when "10111110111",
      "11011101001110001101000000001001100110110111110010011100001111001010100000010111110100010011100000111101" when "10111111000",
      "11011101001110001101000000001001100110110111110010011100001111001010100000010111110100010011100000111101" when "10111111001",
      "11011101010101001100000011111001110000010010010111110110010000010000000011101100111101010001101111000001" when "10111111010",
      "11011101011100001011010011110110111100010111101001100111001011101011101111110110000011100010110000001000" when "10111111011",
      "11011101011100001011010011110110111100010111101001100111001011101011101111110110000011100010110000001000" when "10111111100",
      "11011101100011001010110000000001110101110001110110011100100001111011010111101110110100000111000111010110" when "10111111101",
      "11011101101010001010011000011011000111001110101100110101101101011110110000111111010111110000010000110110" when "10111111110",
      "11011101101010001010011000011011000111001110101100110101101101011110110000111111010111110000010000110110" when "10111111111",
      "11011101110001001010001101000011011011011111011011011100100000101101011010001010101011010101001010011100" when "11000000000",
      "11011101111000001010001101111011011101011000110001011101100111000010000110011100101100011000001110010010" when "11000000001",
      "11011101111000001010001101111011011101011000110001011101100111000010000110011100101100011000001110010010" when "11000000010",
      "11011101111111001010011011000011110111110010111111000001001001011101010010000001010101100110010010111011" when "11000000011",
      "11011110000110001010110100011101010101101001110101100011010110011110100010010011110101101100011000011001" when "11000000100",
      "11011110000110001010110100011101010101101001110101100011010110011110100010010011110101101100011000011001" when "11000000101",
      "11011110001101001011011010001000100001111100101000001101001101010101110101011100111011010101110110010111" when "11000000110",
      "11011110001101001011011010001000100001111100101000001101001101010101110101011100111011010101110110010111" when "11000000111",
      "11011110010100001100001100000110000111101110001100001101001100101101000100011101000010110111111001111011" when "11000001000",
      "11011110011011001101001010010110110010000100111001010000000100101010011011100110100101100001000011100010" when "11000001001",
      "11011110011011001101001010010110110010000100111001010000000100101010011011100110100101100001000011100010" when "11000001010",
      "11011110100010001110010100111011001100001010101001111001101100001100001100110010111110110100110100010100" when "11000001011",
      "11011110101001001111101011110100000001001100111011111101111001111110011111100100010011001101001110100110" when "11000001100",
      "11011110101001001111101011110100000001001100111011111101111001111110011111100100010011001101001110100110" when "11000001101",
      "11011110110000010001001111000001111100011100110000111001100000101011100010101011111010001101001111010010" when "11000001110",
      "11011110110111010010111110100101101001001110101110001011001110100111000011010101101000100001001011111001" when "11000001111",
      "11011110110111010010111110100101101001001110101110001011001110100111000011010101101000100001001011111001" when "11000010000",
      "11011110111110010100111010011111110010111010111101101100110000110101001101111101110000011101100011101110" when "11000010001",
      "11011111000101010111000010110001000100111101001110001011111001101101111100111111001100000000101010110111" when "11000010010",
      "11011111000101010111000010110001000100111101001110001011111001101101111100111111001100000000101010110111" when "11000010011",
      "11011111001100011001010111011010001010110100110011100011101010111100111001101110000001010001111001101110" when "11000010100",
      "11011111010011011011111000011011110000000100100111010101100010111110110011111001110001110001010100101111" when "11000010101",
      "11011111010011011011111000011011110000000100100111010101100010111110110011111001110001110001010100101111" when "11000010110",
      "11011111011010011110100101110110100000010011001001000010101101111100110100011001100101100101000111000010" when "11000010111",
      "11011111011010011110100101110110100000010011001001000010101101111100110100011001100101100101000111000010" when "11000011000",
      "11011111100001100001011111101011000111001010011110100101011010000110001111101011100110001111100101110000" when "11000011001",
      "11011111101000100100100101111010010000011000010100101010001111101001011100111000000000111001011100100110" when "11000011010",
      "11011111101000100100100101111010010000011000010100101010001111101001011100111000000000111001011100100110" when "11000011011",
      "11011111101111100111111000100100100111101101111111001001101100001100010110001111001100111111110100010001" when "11000011100",
      "11011111110110101011010111101010111001000000011001100001100001100101001000000001011011111110010011100100" when "11000011101",
      "11011111110110101011010111101010111001000000011001100001100001100101001000000001011011111110010011100100" when "11000011110",
      "11011111111101101111000011001101110000001000000111001110011000010011110010110101111110111001100011110111" when "11000011111",
      "11100000000100110010111011001101111001000001010100000101010101011101000110101110011001100000011011001110" when "11000100000",
      "11100000000100110010111011001101111001000001010100000101010101011101000110101110011001100000011011001110" when "11000100001",
      "11100000001011110110111111101011111111101011110100101101100100000111011100001010000101110000010001000100" when "11000100010",
      "11100000010010111011010000101000110000001011000110111010000010011010010000100101011000100101001001100000" when "11000100011",
      "11100000010010111011010000101000110000001011000110111010000010011010010000100101011000100101001001100000" when "11000100100",
      "11100000011001111111101110000100110110100110010010000011010010000000101011110110100111100000100101101100" when "11000100101",
      "11100000011001111111101110000100110110100110010010000011010010000000101011110110100111100000100101101100" when "11000100110",
      "11100000100001000100011000000000111111001000000111100001001100001111110100010010111111011010000000101111" when "11000100111",
      "11100000101000001001001110011101110101111111000011000100111001110001010111001100001110111011001000101011" when "11000101000",
      "11100000101000001001001110011101110101111111000011000100111001110001010111001100001110111011001000101011" when "11000101001",
      "11100000101111001110010001011100000111011101001011010010101101110011001011011111011011000000110011100100" when "11000101010",
      "11100000110110010011100000111100011111111000010001111100000100111100010100110100101001010110100100100111" when "11000101011",
      "11100000110110010011100000111100011111111000010001111100000100111100010100110100101001010110100100100111" when "11000101100",
      "11100000111101011000111100111111101011101001110100011001100111101000001100110110100011101001000100010101" when "11000101101",
      "11100001000100011110100101100110010111001110111100000101010000001000011001010000001111011001010101001100" when "11000101110",
      "11100001000100011110100101100110010111001110111100000101010000001000011001010000001111011001010101001100" when "11000101111",
      "11100001001011100100011010110001001111001000011110110100010100001101110100100111010000010010000011110111" when "11000110000",
      "11100001001011100100011010110001001111001000011110110100010100001101110100100111010000010010000011110111" when "11000110001",
      "11100001010010101010011100100000111111111010111111010001110010011001110000101111000110111111110010101101" when "11000110010",
      "11100001011001110000101010110110010110001110101101011000100010110111011000111010111100010110100101011010" when "11000110011",
      "11100001011001110000101010110110010110001110101101011000100010110111011000111010111100010110100101011010" when "11000110100",
      "11100001100000110111000101110001111110101111100110101101101011111110011010111001100111100011010101010001" when "11000110101",
      "11100001100111111101101101010100100110001101010110111010111010011111011101001111111111100100110100010100" when "11000110110",
      "11100001100111111101101101010100100110001101010110111010111010011111011101001111111111100100110100010100" when "11000110111",
      "11100001101111000100100001011110111001011011011000001000111101011010101010001100101010010001010110011010" when "11000111000",
      "11100001110110001011100010010001100101010000110011011010000101100001010101111000000000000001111000000001" when "11000111001",
      "11100001110110001011100010010001100101010000110011011010000101100001010101111000000000000001111000000001" when "11000111010",
      "11100001111101010010101111101101010110101000100001000100101000100011000111001011000000111011000011011011" when "11000111011",
      "11100001111101010010101111101101010110101000100001000100101000100011000111001011000000111011000011011011" when "11000111100",
      "11100010000100011010001001110010111010100001001001001101101000000111001010011110111111111000100011001100" when "11000111101",
      "11100010001011100001110000100010111101111101000100000011011100010010010101101111110001110110111110011010" when "11000111110",
      "11100010001011100001110000100010111101111101000100000011011100010010010101101111110001110110111110011010" when "11000111111",
      "11100010010010101001100011111110001110000010011010011000100001111010100101010001111001111110000010110101" when "11001000000",
      "11100010011001110001100100000101010111111011000101111110001100101000011001000101111000011110111111011110" when "11001000001",
      "11100010011001110001100100000101010111111011000101111110001100101000011001000101111000011110111111011110" when "11001000010",
      "11100010100000111001110000111001001000110100110001111111011100100110111010011001010000111011100001000101" when "11001000011",
      "11100010101000000010001010011010001110000000111011011011111000000011010001001110001011110111111110011101" when "11001000100",
      "11100010101000000010001010011010001110000000111011011011111000000011010001001110001011110111111110011101" when "11001000101",
      "11100010101111001010110000101001010100110100110001100010101000011011110010001001101010111000100110111100" when "11001000110",
      "11100010101111001010110000101001010100110100110001100010101000011011110010001001101010111000100110111100" when "11001000111",
      "11100010110110010011100011100111001010101001010110001101011011011111101100010000111000110101101110001111" when "11001001000",
      "11100010111101011100100011010100011100111011011110011011100111111111111111100101010110001110011001111110" when "11001001001",
      "11100010111101011100100011010100011100111011011110011011100111111111111111100101010110001110011001111110" when "11001001010",
      "11100011000100100101101111110001111001001011110010101101010110010010000100010111111000001100111010010000" when "11001001011",
      "11100011001011101111001001000000001100111110101111011110101100100100101011110010001010001011110011110110" when "11001001100",
      "11100011001011101111001001000000001100111110101111011110101100100100101011110010001010001011110011110110" when "11001001101",
      "11100011010010111000101111000000000101111100100101100010111111001000000010011110011100010111110100110011" when "11001001110",
      "11100011010010111000101111000000000101111100100101100010111111001000000010011110011100010111110100110011" when "11001001111",
      "11100011011010000010100001110010010001110001011010100000000100001001011101111101000110001000001110011101" when "11001010000",
      "11100011100001001100100001010111011110001101001001001001101011100011011101011111100001010111100000100000" when "11001010001",
      "11100011100001001100100001010111011110001101001001001001101011100011011101011111100001010111100000100000" when "11001010010",
      "11100011101000010110101101110000011001000011100001111100111010100010100111101000000100000111111010011110" when "11001010011",
      "11100011101111100001000110111101110000001100001011011011101011000000001101010110011111010011111001111010" when "11001010100",
      "11100011101111100001000110111101110000001100001011011011101011000000001101010110011111010011111001111010" when "11001010101",
      "11100011110110101011101101000000010001100010100010101000001110110010111100010000101101010010001111110101" when "11001010110",
      "11100011110110101011101101000000010001100010100010101000001110110010111100010000101101010010001111110101" when "11001010111",
      "11100011111101110110011111111000101011000101111011100000110110110110101000111111100000010000011101011011" when "11001011000",
      "11100100000101000001011111100111101010111001100001011011011110001011011011011111000111110101011010000101" when "11001011001",
      "11100100000101000001011111100111101010111001100001011011011110001011011011011111000111110101011010000101" when "11001011010",
      "11100100001100001100101100001101111111000100010111100001011000101101000110101011101110000001010011001000" when "11001011011",
      "11100100010011011000000101101100010101110001011001001011000110000011010101011001110110111000101011010101" when "11001011100",
      "11100100010011011000000101101100010101110001011001001011000110000011010101011001110110111000101011010101" when "11001011101",
      "11100100011010100011101100000011011101001111011010011100001000001011010110010011011010110101101100010001" when "11001011110",
      "11100100011010100011101100000011011101001111011010011100001000001011010110010011011010110101101100010001" when "11001011111",
      "11100100100001101111011111010100000011110001001000011110111101111011110000111001100001111110011011000001" when "11001100000",
      "11100100101000111011011111011110110111101101001010000001000001100011001101110100010111011000110010100100" when "11001100001",
      "11100100101000111011011111011110110111101101001010000001000001100011001101110100010111011000110010100100" when "11001100010",
      "11100100110000000111101100100100100111011101111111101110101011000010011100100001111101100101000101100101" when "11001100011",
      "11100100110000000111101100100100100111011101111111101110101011000010011100100001111101100101000101100101" when "11001100100",
      "11100100110111010100000110100110000001100010000100101111010110100010100000111101100001001111110111000100" when "11001100101",
      "11100100111110100000101101100011110100011011101111000001101110100111110011100000111101101011010000110110" when "11001100110",
      "11100100111110100000101101100011110100011011101111000001101110100111110011100000111101101011010000110110" when "11001100111",
      "11100101000101101101100001011110101110110001001111110111111010100010011110001010111101110111100001110111" when "11001101000",
      "11100101001100111010100010010111011111001100110100010011110000011101000001011011111111010010010111100100" when "11001101001",
      "11100101001100111010100010010111011111001100110100010011110000011101000001011011111111010010010111100100" when "11001101010",
      "11100101010100000111110000001110110100011100100101100011001011101001101100000101010110101110010110110110" when "11001101011",
      "11100101010100000111110000001110110100011100100101100011001011101001101100000101010110101110010110110110" when "11001101100",
      "11100101011011010101001011000101011101010010101001011100100110101111010000101101110101010110001111000101" when "11001101101",
      "11100101100010100010110010111100001000100101000010111011011001110110000100010111101011011100111011111000" when "11001101110",
      "11100101100010100010110010111100001000100101000010111011011001110110000100010111101011011100111011111000" when "11001101111",
      "11100101101001110000100111110011100101001101110010011100011100110101110001011100100111110010100111100110" when "11001110000",
      "11100101101001110000100111110011100101001101110010011100011100110101110001011100100111110010100111100110" when "11001110001",
      "11100101110000111110101001101100100010001010110110011010101101100100101010011100110101101001100000100101" when "11001110010",
      "11100101111000001100111000100111101110011110001011101011111010001001001000000110100001000011010011101000" when "11001110011",
      "11100101111000001100111000100111101110011110001011101011111010001001001000000110100001000011010011101000" when "11001110100",
      "11100101111111011011010100100101111001001101101101111101001111001101111110100100001111101010000000101011" when "11001110101",
      "11100110000110101001111101100111110001100011011000010000001010011010010101101001000101111101100000100101" when "11001110110",
      "11100110000110101001111101100111110001100011011000010000001010011010010101101001000101111101100000100101" when "11001110111",
      "11100110001101111000110011101110000110101101000101010111010000101101101111111001111011100010110101101101" when "11001111000",
      "11100110001101111000110011101110000110101101000101010111010000101101101111111001111011100010110101101101" when "11001111001",
      "11100110010101000111110110111001100111111100110000010011001001000001001100111100001110000011000010011101" when "11001111010",
      "11100110011100010111000111001011000100101000010100101111011010101101110010111011010001100110100011100111" when "11001111011",
      "11100110011100010111000111001011000100101000010100101111011010101101110010111011010001100110100011100111" when "11001111100",
      "11100110100011100110100100100011001100001001101111011111110000011001101011111101101110010111101101011100" when "11001111101",
      "11100110100011100110100100100011001100001001101111011111110000011001101011111101101110010111101101011100" when "11001111110",
      "11100110101010110110001111000010101101111110111110111100111110101100000011101101101101110011001100101110" when "11001111111",
      "11100110110010000110000110101010011001101010000011100010001111001000110001111111001111001001101110110010" when "11010000000",
      "11100110110010000110000110101010011001101010000011100010001111001000110001111111001111001001101110110010" when "11010000001",
      "11100110111001010110001011011010111110110001000000001010001111010100011111001000110001110001110111000000" when "11010000010",
      "11100110111001010110001011011010111110110001000000001010001111010100011111001000110001110001110111000000" when "11010000011",
      "11100111000000100110011101010101001100111101111010101100100100000001101111001011011100100101101100100100" when "11010000100",
      "11100111000111110110111100011001110011111110111100011011000000101000000000110000100101000101110010110100" when "11010000101",
      "11100111000111110110111100011001110011111110111100011011000000101000000000110000100101000101110010110100" when "11010000110",
      "11100111001111000111101000101001100011100110010010011111000010100101001101001011110101011001101000010010" when "11010000111",
      "11100111001111000111101000101001100011100110010010011111000010100101001101001011110101011001101000010010" when "11010001000",
      "11100111010110011000100010000101001011101010001110010111010001001010010110111001101111100111010111101001" when "11010001001",
      "11100111011101101001101000101101011100000101000110010101000001010100010011111011101110000000011001111100" when "11010001010",
      "11100111011101101001101000101101011100000101000110010101000001010100010011111011101110000000011001111100" when "11010001011",
      "11100111100100111010111100100011000100110101010101111001111101110001000001111011100010100111000100110110" when "11010001100",
      "11100111101100001100011101100110110101111101011110010101110011010010010001101001011101111100100011011100" when "11010001101",
      "11100111101100001100011101100110110101111101011110010101110011010010010001101001011101111100100011011100" when "11010001110",
      "11100111110011011110001011111001011111100100000111000100000001001110010111110001001011110100100110000111" when "11010001111",
      "11100111110011011110001011111001011111100100000111000100000001001110010111110001001011110100100110000111" when "11010010000",
      "11100111111010110000000111011011110001110011111110001001101110001111110001001010111110100000010000000111" when "11010010001",
      "11101000000010000010010000001110011100111011111000110011100001010100001000110111101011111001010001100000" when "11010010010",
      "11101000000010000010010000001110011100111011111000110011100001010100001000110111101011111001010001100000" when "11010010011",
      "11101000001001010100100110010010010001001110110011110011011110111011101101111111001101110110010100000101" when "11010010100",
      "11101000001001010100100110010010010001001110110011110011011110111011101101111111001101110110010100000101" when "11010010101",
      "11101000010000100111001001100111111111000011110011111111001010101001101000010010100110010100101100110001" when "11010010110",
      "11101000010111111001111010010000010110110110000110101101101100110101111001111011111001110000000010000011" when "11010010111",
      "11101000010111111001111010010000010110110110000110101101101100110101111001111011111001110000000010000011" when "11010011000",
      "11101000011111001100111000001100001001000101000010010101111100110001111101001111100101110010101110110110" when "11010011001",
      "11101000011111001100111000001100001001000101000010010101111100110001111101001111100101110010101110110110" when "11010011010",
      "11101000100110100000000011011100000110010100000110101100101111000000001101011100010000100101011010011011" when "11010011011",
      "11101000101101110011011100000000111111001010111101100011000111111111101001011111000100100110001011100001" when "11010011100",
      "11101000101101110011011100000000111111001010111101100011000111111111101001011111000100100110001011100001" when "11010011101",
      "11101000110101000111000001111011100100010101011011000100110011001100000000001100100111011101001011001001" when "11010011110",
      "11101000110101000111000001111011100100010101011011000100110011001100000000001100100111011101001011001001" when "11010011111",
      "11101000111100011010110101001100100110100011011110010110011110010011010101000111010110011001011101000100" when "11010100000",
      "11101001000011101110110101110100110110101001010001110100011001000001101101100110010001100001001011100110" when "11010100001",
      "11101001000011101110110101110100110110101001010001110100011001000001101101100110010001100001001011100110" when "11010100010",
      "11101001001011000011000011110101000101011111001011110000111001000011110101110111111111101010100110111100" when "11010100011",
      "11101001001011000011000011110101000101011111001011110000111001000011110101110111111111101010100110111100" when "11010100100",
      "11101001010010010111011111001110000100000001101110110011000010100001001101110111110111101001001000000100" when "11010100101",
      "11101001011001101100001000000000100011010001101010010101010100101110101101110100100000011011001001010011" when "11010100110",
      "11101001011001101100001000000000100011010001101010010101010100101110101101110100100000011011001001010011" when "11010100111",
      "11101001100001000000111110001101010100010011111011000100011011011010010010110000100001010011011101110000" when "11010101000",
      "11101001100001000000111110001101010100010011111011000100011011011010010010110000100001010011011101110000" when "11010101001",
      "11101001101000010110000001110101001000010001101011011110000100010000100011010000000100010011100010100001" when "11010101010",
      "11101001101111101011010010111000110000011000010100001111111000111100111100101111011000110100010011111010" when "11010101011",
      "11101001101111101011010010111000110000011000010100001111111000111100111100101111011000110100010011111010" when "11010101100",
      "11101001110111000000110001011000111101111001011100110110011101100101011010001000010010010001100011000001" when "11010101101",
      "11101001110111000000110001011000111101111001011100110110011101100101011010001000010010010001100011000001" when "11010101110",
      "11101001111110010110011101010110100010001010111011111100010011100010000100010110001110110000100001101110" when "11010101111",
      "11101001111110010110011101010110100010001010111011111100010011100010000100010110001110110000100001101110" when "11010110000",
      "11101010000101101100010110110010001110100110110111111001000000110001111101110010100011101111000000011111" when "11010110001",
      "11101010001101000010011101101100110100101011100111010000011011101101011001101100000011101011010000100010" when "11010110010",
      "11101010001101000010011101101100110100101011100111010000011011101101011001101100000011101011010000100010" when "11010110011",
      "11101010010100011000110010000111000101111011110001010001111011010110110000100111000110001010001001001011" when "11010110100",
      "11101010010100011000110010000111000101111011110001010001111011010110110000100111000110001010001001001011" when "11010110101",
      "11101010011011101111010100000001110011111110001110010111101100001010100011011101010101000101011000100101" when "11010110110",
      "11101010100011000110000011011101110000011110001000100110001001001111011110011101111101000010110000110000" when "11010110111",
      "11101010100011000110000011011101110000011110001000100110001001001111011110011101111101000010110000110000" when "11010111000",
      "11101010101010011101000000011011101101001010111100001011011010000111001101111001011100011101110010101000" when "11010111001",
      "11101010101010011101000000011011101101001010111100001011011010000111001101111001011100011101110010101000" when "11010111010",
      "11101010110001110100001010111100011011111000010111111110110101000000110110001101101101001000110101011001" when "11010111011",
      "11101010111001001011100011000000101110011110011110000000100101101101100001110001100101111001010111010000" when "11010111100",
      "11101010111001001011100011000000101110011110011110000000100101101101100001110001100101111001010111010000" when "11010111101",
      "11101011000000100011001000101001010110111001100011111001011000111000010110001000110110110101101101001111" when "11010111110",
      "11101011000000100011001000101001010110111001100011111001011000111000010110001000110110110101101101001111" when "11010111111",
      "11101011000111111010111011110111000111001010010011011010001100000010000011010011101001010001101101101111" when "11011000000",
      "11101011001111010010111100101010110001010101101010111100000010000001011111010110110101110011111110001010" when "11011000001",
      "11101011001111010010111100101010110001010101101010111100000010000001011111010110110101110011111110001010" when "11011000010",
      "11101011010110101011001011000101000111100100111101111111111100001001100001000100101110011111000100010101" when "11011000011",
      "11101011010110101011001011000101000111100100111101111111111100001001100001000100101110011111000100010101" when "11011000100",
      "11101011011110000011100111000110111100000101110101101110110111110101001100010111101000110010100111011001" when "11011000101",
      "11101011011110000011100111000110111100000101110101101110110111110101001100010111101000110010100111011001" when "11011000110",
      "11101011100101011100010000110001000001001010010001011001110000111011000011011010100011100110110001101000" when "11011000111",
      "11101011101100110101001000000100001001001000100110111001101000101000001111100101110111101011101011000010" when "11011001000",
      "11101011101100110101001000000100001001001000100110111001101000101000001111100101110111101011101011000010" when "11011001001",
      "11101011110100001110001101000001000110011011100011001111110001000100010101100000110110010100110011010010" when "11011001010",
      "11101011110100001110001101000001000110011011100011001111110001000100010101100000110110010100110011010010" when "11011001011",
      "11101011111011100111011111101000101011100010001011000101111101011110100111100010110001010000000001101000" when "11011001100",
      "11101100000011000000111111111011101010111111111011001110110111000101101010011001000000011000100111011010" when "11011001101",
      "11101100000011000000111111111011101010111111111011001110110111000101101010011001000000011000100111011010" when "11011001110",
      "11101100001010011010101101111010110111011100101001000110010110101001111111100001110110100001101001110101" when "11011001111",
      "11101100001010011010101101111010110111011100101001000110010110101001111111100001110110100001101001110101" when "11011010000",
      "11101100010001110100101001100111000011100100100011010010000010101100101001010110010100011000100101001100" when "11011010001",
      "11101100010001110100101001100111000011100100100011010010000010101100101001010110010100011000100101001100" when "11011010010",
      "11101100011001001110110011000001000010001000010010000001110010011010011101000111101010100001011011101100" when "11011010011",
      "11101100100000101001001010001001100101111100110111110000010101010100110110111111111110001010111000011011" when "11011010100",
      "11101100100000101001001010001001100101111100110111110000010101010100110110111111111110001010111000011011" when "11011010101",
      "11101100101000000011101111000001100001111011110001100011111111101001000100011111101010110001011000100011" when "11011010110",
      "11101100101000000011101111000001100001111011110001100011111111101001000100011111101010110001011000100011" when "11011010111",
      "11101100101111011110100001101001101001000010110111101111011011010110011001111100100010011110111110110011" when "11011011000",
      "11101100110110111001100010000010101110010100011110010010011110000100100111110001011010101001011011100011" when "11011011001",
      "11101100110110111001100010000010101110010100011110010010011110000100100111110001011010101001011011100011" when "11011011010",
      "11101100111110010100110000001101100100110111010101011011000011101011000100011000011110100010110101100110" when "11011011011",
      "11101100111110010100110000001101100100110111010101011011000011101011000100011000011110100010110101100110" when "11011011100",
      "11101101000101110000001100001010111111110110101010000110001101101001011111110100110010100010100111001101" when "11011011101",
      "11101101000101110000001100001010111111110110101010000110001101101001011111110100110010100010100111001101" when "11011011110",
      "11101101001101001011110101111011110010100010000110100001000111010011010110011010100011111101111010001011" when "11011011111",
      "11101101010100100111101101100000110000001101110010101010001110101110010111110000010110111000011100111001" when "11011100000",
      "11101101010100100111101101100000110000001101110010101010001110101110010111110000010110111000011100111001" when "11011100001",
      "11101101011100000011110010111010101100010010010100110010100010100101010111101110011010001001011101101110" when "11011100010",
      "11101101011100000011110010111010101100010010010100110010100010100101010111101110011010001001011101101110" when "11011100011",
      "11101101100011100000000110001010011010001100110001111110110100101111111111001100000100000100111000110010" when "11011100100",
      "11101101100011100000000110001010011010001100110001111110110100101111111111001100000100000100111000110010" when "11011100101",
      "11101101101010111100100111010000101101011110101110101001000001110000010010010110010110001111111100010011" when "11011100110",
      "11101101110010011001010110001110011001101110001111000001101101000111000010110101100110000001111111100101" when "11011100111",
      "11101101110010011001010110001110011001101110001111000001101101000111000010110101100110000001111111100101" when "11011101000",
      "11101101111001110110010011000100010010100101110111110001100010011111100011110011001000110000001110110011" when "11011101001",
      "11101101111001110110010011000100010010100101110111110001100010011111100011110011001000110000001110110011" when "11011101010",
      "11101110000001010011011101110011001011110100101110011010111011110011110110011011000110100100101010101100" when "11011101011",
      "11101110001000110000110110011011111001001110011001111011101100001010000101100001011101100111111010100100" when "11011101100",
      "11101110001000110000110110011011111001001110011001111011101100001010000101100001011101100111111010100100" when "11011101101",
      "11101110010000001110011100111111001110101011000011001110101111101100000110111100101000010001111100100111" when "11011101110",
      "11101110010000001110011100111111001110101011000011001110101111101100000110111100101000010001111100100111" when "11011101111",
      "11101110010111101100010001011110000000000111010101101110000000011001111001110011000101001001000111110010" when "11011110000",
      "11101110010111101100010001011110000000000111010101101110000000011001111001110011000101001001000111110010" when "11011110001",
      "11101110011111001010010011111001000001100100011111110100001111110111111000100100101101110000111101101101" when "11011110010",
      "11101110100110101000100100010001000111001000010011011111000101111001110110100011111010001100001000101101" when "11011110011",
      "11101110100110101000100100010001000111001000010011011111000101111001110110100011111010001100001000101101" when "11011110100",
      "11101110101110000111000010100111000100111101000110110001000100001011011111111101100010111111011011110101" when "11011110101",
      "11101110101110000111000010100111000100111101000110110001000100001011011111111101100010111111011011110101" when "11011110110",
      "11101110110101100101101110111011101111010001110100010011101110110111010100011010101001110111001101111110" when "11011110111",
      "11101110110101100101101110111011101111010001110100010011101110110111010100011010101001110111001101111110" when "11011111000",
      "11101110111101000100101001001111111010011001111011111001111010001100110011110001101001101110000010101000" when "11011111001",
      "11101111000100100011110001100100011010101101100011000001111101000110110101001000101010111011001110111011" when "11011111010",
      "11101111000100100011110001100100011010101101100011000001111101000110110101001000101010111011001110111011" when "11011111011",
      "11101111001100000011000111111010000100101001010101011000001000110011000000010101110110100011010100000111" when "11011111100",
      "11101111001100000011000111111010000100101001010101011000001000110011000000010101110110100011010100000111" when "11011111101",
      "11101111010011100010101100010001101100101110100101011001000101011011000010010110000100100011010001101000" when "11011111110",
      "11101111010011100010101100010001101100101110100101011001000101011011000010010110000100100011010001101000" when "11011111111",
      "11101111011011000010011110101100000111100011001100110100010011110000110100111110000100011011100001110010" when "11100000000",
      "11101111100010100010011111001010001001110001101101001110110011111110010010110101100110011000011101110101" when "11100000001",
      "11101111100010100010011111001010001001110001101101001110110011111110010010110101100110011000011101110101" when "11100000010",
      "11101111101010000010101101101100101000001001010000100101110001011001110000010111110011111101110100011101" when "11100000011",
      "11101111101010000010101101101100101000001001010000100101110001011001110000010111110011111101110100011101" when "11100000100",
      "11101111110001100011001010010100010111011101101001110001010011011111110010111111110011001111111111011110" when "11100000101",
      "11101111110001100011001010010100010111011101101001110001010011011111110010111111110011001111111111011110" when "11100000110",
      "11101111111001000011110101000010001100100111010101000111010011110011011111110011111101111100000111101010" when "11100000111",
      "11110000000000100100101101110110111100100011011000111110011001000101111011001110100111010101011000111100" when "11100001000",
      "11110000000000100100101101110110111100100011011000111110011001000101111011001110100111010101011000111100" when "11100001001",
      "11110000001000000101110100110011011100010011100110010000110111100101110011001110000000000100111001000000" when "11100001010",
      "11110000001000000101110100110011011100010011100110010000110111100101110011001110000000000100111001000000" when "11100001011",
      "11110000001111100111001001111000100000111110011000111111110110011000001110000001111101100001110000100010" when "11100001100",
      "11110000001111100111001001111000100000111110011000111111110110011000001110000001111101100001110000100010" when "11100001101",
      "11110000010111001000101101000110111111101110111000110110011001111011010111011001000100010010010000100001" when "11100001110",
      "11110000010111001000101101000110111111101110111000110110011001111011010111011001000100010010010000100001" when "11100001111",
      "11110000011110101010011110011111101101110100111001101100110011110100000110011011010001110100100010001010" when "11100010000",
      "11110000100110001100011110000011100000100100111100001011110111100111010110101100000000011111101111010001" when "11100010001",
      "11110000100110001100011110000011100000100100111100001011110111100111010110101100000000011111101111010001" when "11100010010",
      "11110000101101101110101011110011001101011000001110010000010101000000001110111001100011010100111010111100" when "11100010011",
      "11110000101101101110101011110011001101011000001110010000010101000000001110111001100011010100111010111100" when "11100010100",
      "11110000110101010001000111101111101001101100101011101110010111000011110000001011111011110011000110011010" when "11100010101",
      "11110000110101010001000111101111101001101100101011101110010111000011110000001011111011110011000110011010" when "11100010110",
      "11110000111100110011110001111001101011000100111110110101001000110011001000110001010011110100001011111100" when "11100010111",
      "11110001000100010110101010010010000111001000100000110010011110111101100101010010010000100001100011000100" when "11100011000",
      "11110001000100010110101010010010000111001000100000110010011110111101100101010010010000100001100011000100" when "11100011001",
      "11110001001011111001110000111001110011100011011010010110100111000010011100000100100000001111110101010011" when "11100011010",
      "11110001001011111001110000111001110011100011011010010110100111000010011100000100100000001111110101010011" when "11100011011",
      "11110001010011011101000101110001100110000110100100010111111011100100101101111110110110001010111010010101" when "11100011100",
      "11110001010011011101000101110001100110000110100100010111111011100100101101111110110110001010111010010101" when "11100011101",
      "11110001011011000000101000111010010100100111101000010110111101110000111000011101011001101101010000000001" when "11100011110",
      "11110001011011000000101000111010010100100111101000010110111101110000111000011101011001101101010000000001" when "11100011111",
      "11110001100010100100011010010100110101000001000001000010010100010101110100110001100101101010011101010110" when "11100100000",
      "11110001101010001000011010000001111101010001111010111010101111110010000000100101101100011011111001111110" when "11100100001",
      "11110001101010001000011010000001111101010001111010111010101111110010000000100101101100011011111001111110" when "11100100010",
      "11110001110001101100101000000010100011011110010100110111010011110101101100001000010010100001000000011101" when "11100100011",
      "11110001110001101100101000000010100011011110010100110111010011110101101100001000010010100001000000011101" when "11100100100",
      "11110001111001010001000100010111011101101111000000101001100110011011001010100000001111100011101111100100" when "11100100101",
      "11110001111001010001000100010111011101101111000000101001100110011011001010100000001111100011101111100100" when "11100100110",
      "11110010000000110101101111000001100010010001100011100010000011110110000000110110101000001110000011111011" when "11100100111",
      "11110010000000110101101111000001100010010001100011100010000011110110000000110110101000001110000011111011" when "11100101000",
      "11110010001000011010101000000001100111011000010110110100011000011010010001010000010111110110101111000100" when "11100101001",
      "11110010001111111111101111011000100011011010101000011011111111011100011110011110001001000100110110110110" when "11100101010",
      "11110010001111111111101111011000100011011010101000011011111111011100011110011110001001000100110110110110" when "11100101011",
      "11110010010111100101000101000111001100110100011011100000100111101011100101110101100111000001001100000101" when "11100101100",
      "11110010010111100101000101000111001100110100011011100000100111101011100101110101100111000001001100000101" when "11100101101",
      "11110010011111001010101001001110011010000110101000111010111101000101101100110011111111000100111001111110" when "11100101110",
      "11110010011111001010101001001110011010000110101000111010111101000101101100110011111111000100111001111110" when "11100101111",
      "11110010100110110000011011101111000001110110111111111001011000001000011111110110011011101110100111010000" when "11100110000",
      "11110010100110110000011011101111000001110110111111111001011000001000011111110110011011101110100111010000" when "11100110001",
      "11110010101110010110011100101001111010110000000110100100110010011110100000100001110101000001101111011011" when "11100110010",
      "11110010110101111100101011111111111011100001011010100101100001001010000001000000001010010010010011011010" when "11100110011",
      "11110010110101111100101011111111111011100001011010100101100001001010000001000000001010010010010011011010" when "11100110100",
      "11110010111101100011001001110001111010111111010001101000010100001110101011000110110010100000010111111011" when "11100110101",
      "11110010111101100011001001110001111010111111010001101000010100001110101011000110110010100000010111111011" when "11100110110",
      "11110011000101001001110110000000110000000010111010000011011011111010110001100101101110001100010010100110" when "11100110111",
      "11110011000101001001110110000000110000000010111010000011011011111010110001100101101110001100010010100110" when "11100111000",
      "11110011001100110000110000101101010001101010011011011011110011010001001010001101000101010111011000100100" when "11100111001",
      "11110011001100110000110000101101010001101010011011011011110011010001001010001101000101010111011000100100" when "11100111010",
      "11110011010100010111111001111000010110111000110111001010010000010100101111100010111111110101101111101000" when "11100111011",
      "11110011011011111111010001100010110110110110001001000000111001110110101001110001001100001101000010100111" when "11100111100",
      "11110011011011111111010001100010110110110110001001000000111001110110101001110001001100001101000010100111" when "11100111101",
      "11110011100011100110110111101101101000101111000111110000100010100111111101011110110011011011011111100101" when "11100111110",
      "11110011100011100110110111101101101000101111000111110000100010100111111101011110110011011011011111100101" when "11100111111",
      "11110011101011001110101100011001100011110101100101101110001010010000000000011000000011101001101000011001" when "11101000000",
      "11110011101011001110101100011001100011110101100101101110001010010000000000011000000011101001101000011001" when "11101000001",
      "11110011110010110110101111100111011111100000010001011000100011101000010011010010101100011010010010100010" when "11101000010",
      "11110011110010110110101111100111011111100000010001011000100011101000010011010010101100011010010010100010" when "11101000011",
      "11110011111010011111000001011000010011001010110101111110000000111111000001101011011001100111001101101111" when "11101000100",
      "11110100000010000111100001101100110110010101111100000010000101100001000110100101110000011110100011011111" when "11101000101",
      "11110100000010000111100001101100110110010101111100000010000101100001000110100101110000011110100011011111" when "11101000110",
      "11110100001001110000010000100110000000100111001010000011011100101100110111100101101011000111001110100010" when "11101000111",
      "11110100001001110000010000100110000000100111001010000011011100101100110111100101101011000111001110100010" when "11101001000",
      "11110100010001011001001110000100101001101001000101000001110111001110010110000110101011110000100011011011" when "11101001001",
      "11110100010001011001001110000100101001101001000101000001110111001110010110000110101011110000100011011011" when "11101001010",
      "11110100011001000010011010001001101001001011010001000100001101100110001000000011000000011101011110001010" when "11101001011",
      "11110100011001000010011010001001101001001011010001000100001101100110001000000011000000011101011110001010" when "11101001100",
      "11110100100000101011110100110101110111000010010001111110101000011011111000101001110010110101111101110010" when "11101001101",
      "11110100100000101011110100110101110111000010010001111110101000011011111000101001110010110101111101110010" when "11101001110",
      "11110100101000010101011110001010001011000111101011111000101110011101100010110001100101110010111101000001" when "11101001111",
      "11110100101111111111010110000111011101011010000011110011111000001100000110000001101100010010100101001101" when "11101010000",
      "11110100101111111111010110000111011101011010000011110011111000001100000110000001101100010010100101001101" when "11101010001",
      "11110100110111101001011100101110100101111101000000010001101001010111001000011010110001001101101000011111" when "11101010010",
      "11110100110111101001011100101110100101111101000000010001101001010111001000011010110001001101101000011111" when "11101010011",
      "11110100111111010011110010000000011100111001001001111010010000001000000110010100111000000011011000011011" when "11101010100",
      "11110100111111010011110010000000011100111001001001111010010000001000000110010100111000000011011000011011" when "11101010101",
      "11110101000110111110010101111101111010011100001100000011001001111110010010110110110001100000101000101001" when "11101010110",
      "11110101000110111110010101111101111010011100001100000011001001111110010010110110110001100000101000101001" when "11101010111",
      "11110101001110101001001000100111110110111000110101010101101110011100101010111000010101101001110001010111" when "11101011000",
      "11110101001110101001001000100111110110111000110101010101101110011100101010111000010101101001110001010111" when "11101011001",
      "11110101010110010100001001111111001010100110111000010101111111101010011101001111101111000111001110001000" when "11101011010",
      "11110101011101111111011010000100101110000011001100001001100000100111101010110111000000000000111001111101" when "11101011011",
      "11110101011101111111011010000100101110000011001100001001100000100111101010110111000000000000111001111101" when "11101011100",
      "11110101100101101010111000111001011001101111101100111110010001010110100001100101101001111000100101101010" when "11101011101",
      "11110101100101101010111000111001011001101111101100111110010001010110100001100101101001111000100101101010" when "11101011110",
      "11110101101101010110100110011110000110010011011100110001110000111010110101001000000101101101110001100110" when "11101011111",
      "11110101101101010110100110011110000110010011011100110001110000111010110101001000000101101101110001100110" when "11101100000",
      "11110101110101000010100010110011101100011010100011111000000101010000011001001100100000101000101010010000" when "11101100001",
      "11110101110101000010100010110011101100011010100011111000000101010000011001001100100000101000101010010000" when "11101100010",
      "11110101111100101110101101111011000100110110010001100011001000111001100000101011011100010101100011001001" when "11101100011",
      "11110101111100101110101101111011000100110110010001100011001000111001100000101011011100010101100011001001" when "11101100100",
      "11110110000100011011000111110101001000011100111100101001111110100110100101100000000000100000000111000000" when "11101100101",
      "11110110000100011011000111110101001000011100111100101001111110100110100101100000000000100000000111000000" when "11101100110",
      "11110110001100000111110000100010110000001010000100010000001010110111111101010010011011111110101010100011" when "11101100111",
      "11110110010011110100101000000100110100111110010000001101010011011010111111000101101001011010011011010001" when "11101101000",
      "11110110010011110100101000000100110100111110010000001101010011011010111111000101101001011010011011010001" when "11101101001",
      "11110110011011100001101110011100001111111111010001110100100100100011011110100111000011011011000001101011" when "11101101010",
      "11110110011011100001101110011100001111111111010001110100100100100011011110100111000011011011000001101011" when "11101101011",
      "11110110100011001111000011101001111010011000000100011100011100100010100001101110010000010010111010010000" when "11101101100",
      "11110110100011001111000011101001111010011000000100011100011100100010100001101110010000010010111010010000" when "11101101101",
      "11110110101010111100100111101110101101011000101110000110011100111011110101001000101100011111111100001101" when "11101101110",
      "11110110101010111100100111101110101101011000101110000110011100111011110101001000101100011111111100001101" when "11101101111",
      "11110110110010101010011010101011100010010110100000000111000001111010100101011011111110001001000000111110" when "11101110000",
      "11110110110010101010011010101011100010010110100000000111000001111010100101011011111110001001000000111110" when "11101110001",
      "11110110111010011000011100100001010010101011110111101101011111100111000001111000000001110111011100010000" when "11101110010",
      "11110110111010011000011100100001010010101011110111101101011111100111000001111000000001110111011100010000" when "11101110011",
      "11110111000010000110101101010000110111111000011110101100000101011101101110100001001011100010010001000101" when "11101110100",
      "11110111001001110101001100111011001011100001001100000000000111101001101011101000100010011011101011000100" when "11101110101",
      "11110111001001110101001100111011001011100001001100000000000111101001101011101000100010011011101011000100" when "11101110110",
      "11110111010001100011111011100001000111010000000100011010001110100010011000011000010001101101110110000000" when "11101110111",
      "11110111010001100011111011100001000111010000000100011010001110100010011000011000010001101101110110000000" when "11101111000",
      "11110111011001010010111001000011100100110100011011000110101100001110110111000111111010010110011011000010" when "11101111001",
      "11110111011001010010111001000011100100110100011011000110101100001110110111000111111010010110011011000010" when "11101111010",
      "11110111100001000010000101100011011110000010110010010101111000001110111001111011101011110110101101001000" when "11101111011",
      "11110111100001000010000101100011011110000010110010010101111000001110111001111011101011110110101101001000" when "11101111100",
      "11110111101000110001100001000001101100110100111100000100110001001011011110000001000100111100000101100100" when "11101111101",
      "11110111101000110001100001000001101100110100111100000100110001001011011110000001000100111100000101100100" when "11101111110",
      "11110111110000100001001011011111001011001001111010100101100100101111011101001001011100011000111100010110" when "11101111111",
      "11110111110000100001001011011111001011001001111010100101100100101111011101001001011100011000111100010110" when "11110000000",
      "11110111111000010001000100111100110011000110000001001000011101101001111100010010110101100011000101010000" when "11110000001",
      "11111000000000000001001101011011011110110010110100100100010111111010111110111110001010010011001001110110" when "11110000010",
      "11111000000000000001001101011011011110110010110100100100010111111010111110111110001010010011001001110110" when "11110000011",
      "11111000000111110001100100111100001000011111001011111111111011001100000111000000111110110000111000010001" when "11110000100",
      "11111000000111110001100100111100001000011111001011111111111011001100000111000000111110110000111000010001" when "11110000101",
      "11111000001111100010001011011111101010011111010001011010011011010101101000110000100000110011110000111000" when "11110000110",
      "11111000001111100010001011011111101010011111010001011010011011010101101000110000100000110011110000111000" when "11110000111",
      "11111000010111010011000001000110111111001100100010010100111111010001111011110010100111000111111111101010" when "11110001000",
      "11111000010111010011000001000110111111001100100010010100111111010001111011110010100111000111111111101010" when "11110001001",
      "11111000011111000100000101110011000001000101110000011011101101111111110000110000111000111100100011010010" when "11110001010",
      "11111000011111000100000101110011000001000101110000011011101101111111110000110000111000111100100011010010" when "11110001011",
      "11111000100110110101011001100100101010101111000010001111000001110100110100111001100000100011001011110111" when "11110001100",
      "11111000100110110101011001100100101010101111000010001111000001110100110100111001100000100011001011110111" when "11110001101",
      "11111000101110100110111100011100110110110001110011101101000010000001101100001000100111011101110110101011" when "11110001110",
      "11111000101110100110111100011100110110110001110011101101000010000001101100001000100111011101110110101011" when "11110001111",
      "11111000110110011000101110011100011111111100110110111011000010101000001011000100111011111000011110010011" when "11110010000",
      "11111000110110011000101110011100011111111100110110111011000010101000001011000100111011111000011110010011" when "11110010001",
      "11111000111110001010101111100100100001000100010100101111001010100101011010001001100011000010011101101101" when "11110010010",
      "11111001000101111100111111110101110101000001101101011010000000010000101011100110100100100010100111011101" when "11110010011",
      "11111001000101111100111111110101110101000001101101011010000000010000101011100110100100100010100111011101" when "11110010100",
      "11111001001101101111011111010001010110110011111001010000011100010000001110010010000110011010001110010011" when "11110010101",
      "11111001001101101111011111010001010110110011111001010000011100010000001110010010000110011010001110010011" when "11110010110",
      "11111001010101100010001101111000000001011111001001010101100010100101000111010010100001011011011000101011" when "11110010111",
      "11111001010101100010001101111000000001011111001001010101100010100101000111010010100001011011011000101011" when "11110011000",
      "11111001011101010101001011101010110000001101001000000100100010001111011100111011001000111010110100000110" when "11110011001",
      "11111001011101010101001011101010110000001101001000000100100010001111011100111011001000111010110100000110" when "11110011010",
      "11111001100101001000011000101010011110001100111001111010111011001011111101100011111000100000011111101010" when "11110011011",
      "11111001100101001000011000101010011110001100111001111010111011001011111101100011111000100000011111101010" when "11110011100",
      "11111001101100111011110100111000000110110010111110000010101010101100001101010100110101101101001101011100" when "11110011101",
      "11111001101100111011110100111000000110110010111110000010101010101100001101010100110101101101001101011100" when "11110011110",
      "11111001110100101111100000010100100101011001001110111100011110001010100101101110010010010110010000100110" when "11110011111",
      "11111001110100101111100000010100100101011001001110111100011110001010100101101110010010010110010000100110" when "11110100000",
      "11111001111100100011011011000000110101011111000011001010001100011011010010100101111111111101110011101111" when "11110100001",
      "11111001111100100011011011000000110101011111000011001010001100011011010010100101111111111101110011101111" when "11110100010",
      "11111010000100010111100100111101110010101001001101111001010101011011011000000010101011001110001110100101" when "11110100011",
      "11111010000100010111100100111101110010101001001101111001010101011011011000000010101011001110001110100101" when "11110100100",
      "11111010001100001011111110001100011000100001111111101101101000011111001101001110100001011010100111000100" when "11110100101",
      "11111010001100001011111110001100011000100001111111101101101000011111001101001110100001011010100111000100" when "11110100110",
      "11111010010100000000100110101101100010111001000111001011110001000001011000001010010000111111011110011011" when "11110100111",
      "11111010011011110101011110100010001101100011110001100100001001110011010110111010001000110101100100100110" when "11110101000",
      "11111010011011110101011110100010001101100011110001100100001001110011010110111010001000110101100100100110" when "11110101001",
      "11111010100011101010100101101011010100011100101011011101110110110001000010110110110000111110110000100010" when "11110101010",
      "11111010100011101010100101101011010100011100101011011101110110110001000010110110110000111110110000100010" when "11110101011",
      "11111010101011011111111100001001110011100100000001100001100101011000011010111100010010001011010001100011" when "11110101100",
      "11111010101011011111111100001001110011100100000001100001100101011000011010111100010010001011010001100011" when "11110101101",
      "11111010110011010101100001111110100110111111100001000100110011100110100010000010100000101101011011010000" when "11110101110",
      "11111010110011010101100001111110100110111111100001000100110011100110100010000010100000101101011011010000" when "11110101111",
      "11111010111011001011010111001010101010111010011000110100111101011010111110111001100001101011111001011000" when "11110110000",
      "11111010111011001011010111001010101010111010011000110100111101011010111110111001100001101011111001011000" when "11110110001",
      "11111011000011000001011011101110111011100101011001100010110001000011001011010110101001000000101011001111" when "11110110010",
      "11111011000011000001011011101110111011100101011001100010110001000011001011010110101001000000101011001111" when "11110110011",
      "11111011001010110111101111101100010101010110110110101101101001101110100000101110011001010101000101111111" when "11110110100",
      "11111011001010110111101111101100010101010110110110101101101001101110100000101110011001010101000101111111" when "11110110101",
      "11111011010010101110010011000011110100101010100111001111010001001100101111101000111110010011110010000011" when "11110110110",
      "11111011010010101110010011000011110100101010100111001111010001001100101111101000111110010011110010000011" when "11110110111",
      "11111011011010100101000101110110010110000010000110000111000111110111110001101111001100111000101011010100" when "11110111000",
      "11111011011010100101000101110110010110000010000110000111000111110111110001101111001100111000101011010100" when "11110111001",
      "11111011100010011100001000000100110110000100010011000110010011101010000011111111001100011110100101101110" when "11110111010",
      "11111011100010011100001000000100110110000100010011000110010011101010000011111111001100011110100101101110" when "11110111011",
      "11111011101010010011011001110000010001011101110011011011010101100010111000101000100111101010100000111010" when "11110111100",
      "11111011101010010011011001110000010001011101110011011011010101100010111000101000100111101010100000111010" when "11110111101",
      "11111011110010001010111010111001100101000000110010011110000101111001110000000001100010011111110111111110" when "11110111110",
      "11111011110010001010111010111001100101000000110010011110000101111001110000000001100010011111110111111110" when "11110111111",
      "11111011111010000010101011100001101101100101000010011011110111100010000111110101111000011111011111100101" when "11111000000",
      "11111100000001111010101011101001101000000111111101000011100001100000110000100100101100010110010110010001" when "11111000001",
      "11111100000001111010101011101001101000000111111101000011100001100000110000100100101100010110010110010001" when "11111000010",
      "11111100001001110010111011010010010001101100100100010001101111110011111001001111011111110010010011111000" when "11111000011",
      "11111100001001110010111011010010010001101100100100010001101111110011111001001111011111110010010011111000" when "11111000100",
      "11111100010001101011011010011100100111011011100010111101011010101111100001110001011010010011001111101100" when "11111000101",
      "11111100010001101011011010011100100111011011100010111101011010101111100001110001011010010011001111101100" when "11111000110",
      "11111100011001100100001001001001100110100011001101100100000101001111000100100100111010011111001101000111" when "11111000111",
      "11111100011001100100001001001001100110100011001101100100000101001111000100100100111010011111001101000111" when "11111001000",
      "11111100100001011101000111011010001100010111100010110110100001111101101000010000100110100010001111010010" when "11111001001",
      "11111100100001011101000111011010001100010111100010110110100001111101101000010000100110100010001111010010" when "11111001010",
      "11111100101001010110010101001111010110010010001100100101011111010110001010100100101101110110101001000101" when "11111001011",
      "11111100101001010110010101001111010110010010001100100101011111010110001010100100101101110110101001000101" when "11111001100",
      "11111100110001001111110010101010000001110010100000001110011010011100110110000100101111011010100100101101" when "11111001101",
      "11111100110001001111110010101010000001110010100000001110011010011100110110000100101111011010100100101101" when "11111001110",
      "11111100111001001001011111101011001100011101011111101000011000110010110100001001111110010101000001100001" when "11111001111",
      "11111100111001001001011111101011001100011101011111101000011000110010110100001001111110010101000001100001" when "11111010000",
      "11111101000001000011011100010011110011111101111001110001001001000101101101011101101000011111010011111000" when "11111010001",
      "11111101000001000011011100010011110011111101111001110001001001000101101101011101101000011111010011111000" when "11111010010",
      "11111101001000111101101000100100110110000100001011011010001010111100001010111010110001110010110111111001" when "11111010011",
      "11111101001000111101101000100100110110000100001011011010001010111100001010111010110001110010110111111001" when "11111010100",
      "11111101010000111000000100011111010000100110011111110101111101100000101001111010001001011110010010110110" when "11111010101",
      "11111101010000111000000100011111010000100110011111110101111101100000101001111010001001011110010010110110" when "11111010110",
      "11111101011000110010110000000100000001100000110001100101010101001011110110011011110110100001011100010110" when "11111010111",
      "11111101011000110010110000000100000001100000110001100101010101001011110110011011110110100001011100010110" when "11111011000",
      "11111101100000101101101011010100000110110100101011000100111000001111111110010100110100001000101000100010" when "11111011001",
      "11111101100000101101101011010100000110110100101011000100111000001111111110010100110100001000101000100010" when "11111011010",
      "11111101101000101000110110010000011110101001100111011010100010100110010000110111110111010010111101010011" when "11111011011",
      "11111101101000101000110110010000011110101001100111011010100010100110010000110111110111010010111101010011" when "11111011100",
      "11111101110000100100010000111010000111001100110011000011010000011111111110100100011011100001101100101111" when "11111011101",
      "11111101110000100100010000111010000111001100110011000011010000011111111110100100011011100001101100101111" when "11111011110",
      "11111101111000011111111011010001111110110001001100100000110000011100001100110110111101111111001111110001" when "11111011111",
      "11111101111000011111111011010001111110110001001100100000110000011100001100110110111101111111001111110001" when "11111100000",
      "11111110000000011011110101011001000011101111100101000111011100000011110010001001011011111100011011100010" when "11111100001",
      "11111110000000011011110101011001000011101111100101000111011100000011110010001001011011111100011011100010" when "11111100010",
      "11111110001000010111111111010000010100100110100001101100011000001100101110100100011011110100111011111101" when "11111100011",
      "11111110001000010111111111010000010100100110100001101100011000001100101110100100011011110100111011111101" when "11111100100",
      "11111110010000010100011000111000101111111010011011010011011100000110010110010011111110111111101111000001" when "11111100101",
      "11111110010000010100011000111000101111111010011011010011011100000110010110010011111110111111101111000001" when "11111100110",
      "11111110011000010001000010010011010100010101011111111101011111101111100010100101010101101000011110011101" when "11111100111",
      "11111110011000010001000010010011010100010101011111111101011111101111100010100101010101101000011110011101" when "11111101000",
      "11111110100000001101111011100001000000100111110011010110110001011000011110100101101110001011111100010111" when "11111101001",
      "11111110100000001101111011100001000000100111110011010110110001011000011110100101101110001011111100010111" when "11111101010",
      "11111110101000001011000100100010110011100111001111100101010010010001000110001100011110010101000010010010" when "11111101011",
      "11111110101000001011000100100010110011100111001111100101010010010001000110001100011110010101000010010010" when "11111101100",
      "11111110110000001000011101011001101100001111100101110111011010100101101100001101101100100010110110110000" when "11111101101",
      "11111110110000001000011101011001101100001111100101110111011010100101101100001101101100100010110110110000" when "11111101110",
      "11111110111000000110000110000110101001100010011111010010100100101010111110100101001111010100011010101011" when "11111101111",
      "11111110111000000110000110000110101001100010011111010010100100101010111110100101001111010100011010101011" when "11111110000",
      "11111111000000000011111110101010101010100111011101100001111111011010111110111100101001010100101100100110" when "11111110001",
      "11111111000000000011111110101010101010100111011101100001111111011010111110111100101001010100101100100110" when "11111110010",
      "11111111001000000010000111000110101110101011111011100101101000000100000110100001100001001011011100110000" when "11111110011",
      "11111111001000000010000111000110101110101011111011100101101000000100000110100001100001001011011100110000" when "11111110100",
      "11111111010000000000011111011011110101000011001110100001001011001011101100010100101111001101101111110110" when "11111110101",
      "11111111010000000000011111011011110101000011001110100001001011001011101100010100101111001101101111110110" when "11111110110",
      "11111111010111111111000111101010111101000110100110001011001101000101100101001101111100001101111010100100" when "11111110111",
      "11111111010111111111000111101010111101000110100110001011001101000101100101001101111100001101111010100100" when "11111111000",
      "11111111011111111101111111110101000110010101001101111100011001100001110101100001110001011110101011000010" when "11111111001",
      "11111111011111111101111111110101000110010101001101111100011001100001110101100001110001011110101011000010" when "11111111010",
      "11111111100111111101000111111011010000010100001101011110111010110010001100001100100100100010010011101110" when "11111111011",
      "11111111100111111101000111111011010000010100001101011110111010110010001100001100100100100010010011101110" when "11111111100",
      "11111111101111111100011111111110011010101110101001011101111000001000011111110110010111110101110011011011" when "11111111101",
      "11111111101111111100011111111110011010101110101001011101111000001000011111110110010111110101110011011011" when "11111111110",
      "11111111110111111100000111111111100101010101100100010100111011101111100110011000011101010010011101001101" when "11111111111",
      "--------------------------------------------------------------------------------------------------------" when others;
   Y1_c0 <= Y0_c0; -- for the possible blockram register
   Y <= Y1_c0;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable1_Freq300_uid40
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable1_Freq300_uid40 is
    port (clk, ce_2 : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(94 downto 0)   );
end entity;

architecture arch of LogTable1_Freq300_uid40 is
signal Y0_c2 :  std_logic_vector(94 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c2 :  std_logic_vector(94 downto 0);
signal X_c2 :  std_logic_vector(8 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_2 = '1' then
               X_c2 <= X;
            end if;
         end if;
      end process;
   with X_c2  select  Y0_c2 <= 
      "00000000010000000000000000000011111111111111111110101010101010101011001010101010101010011101111" when "000000000",
      "00000000110000000000000000000100000000000000000001010101010101010101110101010101010101100010001" when "000000001",
      "00000001010000000000000000100100000000000000100100000000000000101000100000000000110000100110011" when "000000010",
      "00000001110000000000000001100100000000000010100110101010101111100011001010110100011011101011000" when "000000011",
      "00000010010000000000000011000100000000000111001001010101101000000101110110001001110110110001011" when "000000100",
      "00000010110000000000000101000100000000001111001100000000110011010000100010111000100001111110000" when "000000101",
      "00000011010000000000000111100100000000011011101110101100011101000011010010100001111101011011100" when "000000110",
      "00000011110000000000001010100100000000101101110001011000110100011110000111011101101001011110000" when "000000111",
      "00000100010000000000001110000100000001000110010100000110001011100001000101000101000110100111110" when "000001000",
      "00000100110000000000010010000100000001100110010110110100110111001100001111111111110101101111011" when "000001001",
      "00000101010000000000010110100100000010001110111001100101001111011111101110001111011000000101110" when "000001010",
      "00000101110000000000011011100100000011000000111100010111101111011011100111011011001111011101110" when "000001011",
      "00000110010000000000100001000100000011111101011111001100110101000000000100111100111110010101000" when "000001100",
      "00000110110000000000100111000100000101000101100010000101000001001101010010001100000111111100101" when "000001101",
      "00000111010000000000101101100100000110011010000101000000111000000011011100101010010000100100000" when "000001110",
      "00000111110000000000110100100100000111111100001000000001000000100010110100001110111101100100001" when "000001111",
      "00001000010000000000111100000100001001101100101011000110000100101011101011010011110101101011011" when "000010000",
      "00001000110000000001000100000100001011101100101110010000110001011110010111000000100001001010110" when "000010001",
      "00001001010000000001001100100100001101111101010001100001110110111011001111010110101010000100011" when "000010010",
      "00001001110000000001010101100100010000011111010100111010001000000010101111011101111100011001111" when "000010011",
      "00001010010000000001011111000100010011010011111000011010011010110101010101110000000110011100110" when "000010100",
      "00001010110000000001101001000100010110011011111100000011101000010011100100000100111000111111000" when "000010101",
      "00001011010000000001110011100100011001111000011111110110101100011101111111111110000111100101010" when "000010110",
      "00001011110000000001111110100100011101101010100011110100100110010101010010110011101000111001000" when "000010111",
      "00001100010000000010001010000100100001110011000111111110010111111010001001111111010110111100110" when "000011000",
      "00001100110000000010010110000100100110010011001100010101000110001101010111001001001111100000110" when "000011001",
      "00001101010000000010100010100100101011001011110000111001111001001111110000010011010100011000000" when "000011010",
      "00001101110000000010101111100100110000011101110101101101111100000010010000000101101011101111010" when "000011011",
      "00001110010000000010111101000100110110001010011010110010011100100101110101111010100000100100000" when "000011100",
      "00001110110000000011001011000100111100010010100000001000101011111011100110001010000010111101101" when "000011101",
      "00001111010000000011011001100101000010110111000101110001111110000100101010010110101000100101110" when "000011110",
      "00001111110000000011101000100101001001111001001011101111101010000010010001011000101101000011011" when "000011111",
      "00010000010000000011111000000101010001011001110010000011001001110101101111101010110010010101011" when "000100000",
      "00010000110000000100001000000101011001011001111000101101111010100000011111010101100001001111000" when "000100001",
      "00010001010000000100011000100101100001111010011111110001011100000100000000011011101001110101000" when "000100010",
      "00010001110000000100101001100101101010111100100111001111010001100001111001000110000011111011100" when "000100011",
      "00010010010000000100111011000101110100100001001111001001000000111011110101101111101111100101000" when "000100100",
      "00010010110000000101001101000101111110101001010111100000010011010011101001010001110101100010000" when "000100101",
      "00010011010000000101011111100110001001010110000000010110110100101011001101001111100111110010010" when "000100110",
      "00010011110000000101110010100110010100101000001001101110010100000100100010000010100010000110010" when "000100111",
      "00010100010000000110000110000110100000100000110011101000100011100001101111000110001010100010010" when "000101000",
      "00010100110000000110011010000110101101000000111110000111011000000101000011000100010010000001100" when "000101001",
      "00010101010000000110101110100110111010001001101001001100101001110000110100000000110100111010110" when "000101010",
      "00010101110000000111000011100111000111111011110100111010010011100111011111100101111011100110010" when "000101011",
      "00010110010000000111011001000111010110011000100001010010010011101011101011001111111011000100010" when "000101100",
      "00010110110000000111101111000111100101100000101110010110101011000000000100011001010101100011100" when "000101101",
      "00010111010000001000000101100111110101010101011100001001011101100111100000100110111011001010110" when "000101110",
      "00010111110000001000011100101000000101110111101010101100110010100100111101110011101010100001000" when "000101111",
      "00011000010000001000110100001000010111001000011010000010110011111011100010011100110001011000101" when "000110000",
      "00011000110000001001001100001000101001001000101010001101101110101110011101101101101101011001101" when "000110001",
      "00011001010000001001100100101000111011111001011011001111110011000001000111101100001100101110101" when "000110010",
      "00011001110000001001111101101001001111011011101101001011010011110111000001100100001110110000111" when "000110011",
      "00011010010000001010010111001001100011110000100000000010100111010011110101110100000100110111011" when "000110100",
      "00011010110000001010110001001001111000111000110011111000000110011011011000011000010011000100101" when "000110101",
      "00011011010000001011001011101010001110110101101000101110001101010001100110110111110000110111100" when "000110110",
      "00011011110000001011100110101010100101100111111110100111011010111010101000101111101001111011001" when "000110111",
      "00011100010000001100000010001010111101010000110101100110010001011010101111011111011110111001010" when "000111000",
      "00011100110000001100011110001011010101110001001101101101010101110110010110110101000110001100100" when "000111001",
      "00011101010000001100111010101011101111001010000110111111010000010010000100111000101100110100011" when "000111010",
      "00011101110000001101010111101100001001011100100001011110101011110010101010011000110111001001011" when "000111011",
      "00011110010000001101110101001100100100101001011101001110010110011101000010110110100001110010110" when "000111100",
      "00011110110000001110010011001101000000110001111010010001000001010110010100110001000010011100100" when "000111101",
      "00011111010000001110110001101101011101110110111000101001100000100011110001110010001000101111100" when "000111110",
      "00011111110000001111010000101101111011111001011000011010101011001010110110111001111111001000111" when "000111111",
      "00100000010000001111110000001110011010111010011001100111011011010001001100101011001011110100000" when "001000000",
      "00100000110000010000010000001110111010111010111100010010101101111100100111010110110001100100000" when "001000001",
      "00100001010000010000110000101111011011111100000000011111100011010011000111001000010000101111101" when "001000010",
      "00100001110000010001010001101111111101111110100110010000111110011010111000010001101000001100100" when "001000011",
      "00100010010000010001110011010000100001000011101101101010000101011010010011010111010110001100101" when "001000100",
      "00100010110000010010010101010001000101001100010110101110000001010111111101011100011001011100000" when "001000101",
      "00100011010000010010110111110001101010011001100001011111111110011010101000001110010001111111111" when "001000110",
      "00100011110000010011011010110010010000101100001110000011001011101001010010010001000010010110000" when "001000111",
      "00100100010000010011111110010010111000000101011100011010111011001011000111001011010000010110000" when "001001000",
      "00100100110000010100100010010011100000100110001100101010100010000111011111110010000110010010010" when "001001001",
      "00100101010000010101000110110100001010001111011110110101011000100110000010010101010011111011100" when "001001010",
      "00100101110000010101101011110100110101000010010010111110111001101110100010101011001111100011100" when "001001011",
      "00100110010000010110010001010101100000111111101001001010100011101001000010011100110111000010000" when "001001100",
      "00100110110000010110110111010110001110001000100001011011110111011101110001010001110000111010000" when "001001101",
      "00100111010000010111011101110110111100011101111011110110011001010101001100111100001101100000011" when "001001110",
      "00100111110000011000000100110111101100000000111000011101110000011000000001100101001000000010110" when "001001111",
      "00101000010000011000101100011000011100110010010111010101100110101111001001111000000111110000010" when "001010000",
      "00101000110000011001010100011001001110110011011000100001101001100011101111001111100001000010011" when "001010001",
      "00101001010000011001111100111010000010000100111100000101101000111111001010000000010110100111000" when "001010010",
      "00101001110000011010100101111010110110101000000010000101011000001011000001100110011010101011110" when "001010011",
      "00101010010000011011001111011011101100011101101010100100101101010001001100110000010000001010001" when "001010100",
      "00101010110000011011111001011100100011100110110101100111100001011011110001101011001011110011111" when "001010101",
      "00101011010000011100100011111101011100000100100011010001110000110101000110001111010101100001100" when "001010110",
      "00101011110000011101001110111110010101110111110011100111011010100111110000001011101001100000100" when "001010111",
      "00101100010000011101111010011111010001000001100110101100100000111110100101010001111001100011111" when "001011000",
      "00101100110000011110100110100000001101100010111100100101001001000100101011100010101110010100000" when "001011001",
      "00101101010000011111010011000001001011011100110101010101011011000101011001011001101000100001000" when "001011010",
      "00101101110000100000000000000010001010110000010001000001100010001100010101111001000010010100110" when "001011011",
      "00101110010000100000101101100011001011011110001111101101101100100101011000110110010000100110110" when "001011100",
      "00101110110000100001011011100100001101100111110001011110001011011100101011000101100100010000011" when "001011101",
      "00101111010000100010001010000101010001001101110110010111010010111110100110100110001011100010110" when "001011110",
      "00101111110000100010111001000110010110010001011110011101011010010111110110101110010011011100010" when "001011111",
      "00110000010000100011101000100111011100110011101001110100111011110101011000010111001001000000101" when "001100000",
      "00110000110000100100011000101000100100110101011000100010010100100100011010001000111010110000101" when "001100001",
      "00110001010000100101001001001001101110010111101010101010000100110010011100100110111010000011100" when "001100010",
      "00110001110000100101111010001010111001011011100000010000101111101101010010011011011100100001001" when "001100011",
      "00110010010000100110101011101100000110000001111001011010111011100011000000100011111101011100101" when "001100100",
      "00110010110000100111011101101101010100001011110110001101010001100001111110011100111111010000110" when "001100101",
      "00110011010000101000010000001110100011111010010110101100011101111000110110001110001100111100110" when "001100110",
      "00110011110000101001000011001111110101001110011010111101001111110110100100110110011011100010001" when "001100111",
      "00110100010000101001110110110001001000001001000011000100011001101010011010010111101011100011010" when "001101000",
      "00110100110000101010101010110010011100101011001111000110110000100011111010000011001010100011110" when "001101001",
      "00110101010000101011011111010011110010110101111111001001001100110010111010100101010100101000010" when "001101010",
      "00110101110000101100010100010101001010101010010011010000101001100111100110010001110101111000110" when "001101011",
      "00110110010000101101001001110110100100001001001011100010000101010010011011001111101100000011000" when "001101100",
      "00110110110000101101111111110111111111010011101000000010100001000100001011100101000111111101110" when "001101101",
      "00110111010000101110110110011001011100001010101000110111000001001101111101100011101111001101010" when "001101110",
      "00110111110000101111101101011010111010101111001110000100101101000001001011110100011101101000111" when "001101111",
      "00111000010000110000100100111100011011000010010111110000101110101111100101100011100111000001011" when "001110000",
      "00111000110000110001011100111101111101000101000110000000010011101011001110101100111000100111111" when "001110001",
      "00111001010000110010010101011111100000111000011000111000101100000110100000000111011010110110010" when "001110010",
      "00111001110000110011001110100001000110011101010000011111001011010100000111110001110010111000011" when "001110011",
      "00111010010000110100001000000010101101110100101100111001000111100111001000111110000100010101111" when "001110100",
      "00111010110000110101000010000100010110111111101110001011111010010010111100011101110010111101011" when "001110101",
      "00111011010000110101111100100110000001111111010100011100111111101011010000101110000100010000101" when "001110110",
      "00111011110000110110110111100111101110110100011111110001110111000100001010000011100001010001000" when "001110111",
      "00111100010000110111110011001001011101100000010000010000000010110010000010110110011000001101100" when "001111000",
      "00111100110000111000101111001011001110000011100101111101001000001001101011101110011110010001100" when "001111001",
      "00111101010000111001101011101101000000011111100000111110101111100000001011101111010001010100110" when "001111010",
      "00111101110000111010101000101110110100110101000001011010100100001011000000100011111001101011101" when "001111011",
      "00111110010000111011100110010000101011000101000111010110010100011111111110101011001011111000110" when "001111100",
      "00111110110000111100100100010010100011010000110010110111110001110101010001100011101010100000000" when "001111101",
      "00111111010000111101100010110100011101011001000100000100110000100001011011110111100111111001010" when "001111110",
      "00111111110000111110100001110110011001011110111011000011000111111011010111101001001000000101100" when "001111111",
      "01000000010000111111100001011000010111100011010111111000110010011010010110011110000010100011101" when "010000000",
      "01000000110001000000100001011010010111100111011010101011101101010110000001101100000100000111011" when "010000001",
      "01000001010001000001100001111100011001101100000011100001111001000110011010100100110000101111110" when "010000010",
      "01000001110001000010100010111110011101110010010010100001011001000011111010100001100101011111110" when "010000011",
      "01000010010001000011100100100000100011111011000111110000010011100111010011001111111010010111110" when "010000100",
      "01000010110001000100100110100010101100000111100011010100110010001001101110111101000100001110100" when "010000101",
      "01000011010001000101101001000100110110011000100101010101000001000100110000100010010110101101001" when "010000110",
      "01000011110001000110101100000111000010101111001101110111001111110010010011110001000110001010111" when "010000111",
      "01000100010001000111101111101001010001001100011101000001110000101100101101011110101001101001101" when "010001000",
      "01000100110001001000110011101011100001110001010010111010111001001110101011110000011100110100000" when "010001001",
      "01000101010001001001111000001101110100011110101111101001000001110011010110001000000001111100001" when "010001010",
      "01000101110001001010111101010000001001010101110011010010100101110110001101101111000011111011000" when "010001011",
      "01000110010001001100000010110010100000010111011101111110000011110011001101100011011000010001110" when "010001100",
      "01000110110001001101001000110100111001100100101111110001111101000110101010100011000001001010100" when "010001101",
      "01000111010001001110001111010111010100111110101000110100110110001101010011111000001111011011101" when "010001110",
      "01000111110001001111010110011001110010100110001001001101010110100100010011000101100100101010011" when "010001111",
      "01001000010001010000011101111100010010011100010001000010001000101001001100010001110101010000000" when "010010000",
      "01001000110001010001100101111110110100100010000000011001111001111001111110010100001010011111000" when "010010001",
      "01001001010001010010101110100001011000111000010111011011011010110101000011000000000100101000110" when "010010010",
      "01001001110001010011110111100011111111100000010110001101011110111001001111010001011101000101100" when "010010011",
      "01001010010001010101000001000110101000011010111100110110111100100101110011011000101000011100011" when "010010100",
      "01001010110001010110001011001001010011101001001011011110101101011010011011000110011000101100000" when "010010101",
      "01001011010001010111010101101100000001001100000010001011101101110111001101110111111111010101000" when "010010110",
      "01001011110001011000100000101110110001000100100001000100111101011100101111000011001111100101000" when "010010111",
      "01001100010001011001101100010001100011010011101000010001011110101011111110000010100000100010100" when "010011000",
      "01001100110001011010111000010100010111111010010111111000010111000110010110100000101111011001010" when "010011001",
      "01001101010001011100000100110111001110111001110000000000101111001101110000100101100001101000110" when "010011010",
      "01001101110001011101010001111010001000010010110000110001110010100100100001000001000111010011000" when "010011011",
      "01001110010001011110011111011101000100000110011010010010101111101101011001011000011101001011010" when "010011100",
      "01001110110001011111101101100000000010010101101100101010111000001011101000010001001111000111110" when "010011101",
      "01001111010001100000111100000011000011000001101000000001100000100010111001011101111010010011000" when "010011110",
      "01001111110001100010001011000110000110001011001100011110000000010111010110001001101111011101100" when "010011111",
      "01010000010001100011011010101001001011110011011010000111110010001101100101000100110101010010100" when "010100000",
      "01010000110001100100101010101100010011111011010001000110010011101010101010110000001010101011011" when "010100001",
      "01010001010001100101111011001111011110100011110001100001000101010100001001101001101001000101010" when "010100010",
      "01010001110001100111001100010010101011101101111011011111101010110000000010011000000110110111100" when "010100011",
      "01010010010001101000011101110101111011011010101111001001101010100100110011110111011001101010100" when "010100100",
      "01010010110001101001101111111001001101101011001100100110101110011001011011100100011000110000101" when "010100101",
      "01010011010001101011000010011100100010100000010011111110100010110101010101101000111111011110010" when "010100110",
      "01010011110001101100010101011111111001111011000101011000110111100000011101001000001111100100110" when "010100111",
      "01010100010001101101101001000011010011111100100000111101011111000011001100001010010011101100100" when "010101000",
      "01010100110001101110111101000110110000100101100110110100001111000110011100001000100001110010001" when "010101001",
      "01010101010001110000010001101010001111110111010111000101000000010011100101111001011101100010000" when "010101010",
      "01010101110001110001100110101101110001110010110001110111101110010100100001111100111010110110110" when "010101011",
      "01010110010001110010111100010001010110011000110111010100010111110011101000101000000000011000010" when "010101100",
      "01010110110001110100010010010100111101101010100111100010111110011011110010010001001001111010100" when "010101101",
      "01010111010001110101101000111000100111101001000010101011100110111000010111011100001010111111000" when "010101110",
      "01010111110001110110111111111100010100010101001000110110011000110101010001000110010001010110000" when "010101111",
      "01011000010001111000010111100000000011101111111010001011011110111110111000110010000111100001000" when "010110000",
      "01011000110001111001101111100011110101111010010110110011000111000010001000110011110111010110000" when "010110001",
      "01011001010001111011001000000111101010110101011110110101100001101100011100011101001100100100101" when "010110010",
      "01011001110001111100100001001011100010100010010010011011000010101011110000001001010111011010100" when "010110011",
      "01011010010001111101111010101111011101000001110001101100000000101110100001101001001111001010001" when "010110100",
      "01011010110001111111010100110011011010010100111100110000110101100011110000001111010100110010001" when "010110101",
      "01011011010010000000101111010111011010011100110011110001111101111010111100111011110101100101000" when "010110110",
      "01011011110010000010001010011011011101011010010110110111111001100100001010101000101101110010110" when "010110111",
      "01011100010010000011100101111111100011001110100110001011001011001111111110010101101011010010010" when "010111000",
      "01011100110010000101000010000011101011111010100001110100011000101111011111010100010000001100110" when "010111001",
      "01011101010010000110011110100111110111011111001001111100001010110100010111010011110101101001101" when "010111010",
      "01011101110010000111111011101100000101111101011110101011001101010000110010101101101110011011100" when "010111011",
      "01011110010010001001011001010000010111010110100000001010001110110111100000110001001001101101100" when "010111100",
      "01011110110010001010110111010100101011101011001110100010000001011011110011101111010101110010101" when "010111101",
      "01011111010010001100010101111001000010111100101001111011011001110001100001000111100010110100110" when "010111110",
      "01011111110010001101110100111101011101001011110010011111001111101101000001110011000101100101111" when "010111111",
      "01100000010010001111010100100001111010011001101000010110011110000011010010010001011010010001011" when "011000000",
      "01100000110010010000110100100110011010100111001011101010000010101001110010110100000111001110110" when "011000001",
      "01100001010010010010010101001010111101110101011100100010111110010110100111101010111111110100110" when "011000010",
      "01100001110010010011110110001111100100000101011011001010010101000000011001010000000111001101110" when "011000011",
      "01100010010010010101010111110100001101011000000111101001001101011110010100010011110011001110000" when "011000100",
      "01100010110010010110111001111000111001101110100010001000110001101000001010001000101111001000010" when "011000101",
      "01100011010010011000011100011101101001001001101010110010001110010110010000101111111110100110100" when "011000110",
      "01100011110010011001111111100010011011101010100001101110110011100001100011000101000000100001101" when "011000111",
      "01100100010010011011100011000111010001010010000111000111110100000011100001001001110001111010000" when "011001000",
      "01100100110010011101000111001100001010000001011011000110100101110110010000010010110000110010011" when "011001001",
      "01100101010010011110101011110001000101111001011101110100100001110100011011010010111111001010000" when "011001010",
      "01100101110010100000010000110110000100111011001111011011000011111001010010101000000101111001110" when "011001011",
      "01100110010010100001110110011011000111000111110000000011101011000000101100100110010111101111010" when "011001100",
      "01100110110010100011011100100000001100011111111111110111111001000111000101100100110100001100110" when "011001101",
      "01100111010010100101000011000101010101000100111111000001010011001001100000001001001010100110000" when "011001110",
      "01100111110010100110101010001010100000110111101101101001100001000101100101010011111101000001010" when "011001111",
      "01101000010010101000010001101111101111111001001011111010001101111001100100101100100011010111010" when "011010000",
      "01101000110010101001111001110101000010001010011001111101000111100100010100101101001110010101000" when "011010001",
      "01101001010010101011100010011010010111101100010111111011111111000101010010101111001010011110100" when "011010010",
      "01101001110010101101001011011111110000100000000110000000101000011100100011010110100011010001011" when "011010011",
      "01101010010010101110110101000101001100100110100100010100111010101010110010011110100110001010101" when "011010100",
      "01101010110010110000011111001010101100000000110011000010101111110001010011100101100101101010110" when "011010101",
      "01101011010010110010001001110000001110101111110010010100000100110010000001111000111100011100110" when "011010110",
      "01101011110010110011110100110101110100110100100010010010111001101111100000100001010000011101000" when "011010111",
      "01101100010010110101100000011011011110010000000011001001010001101100111010101110010110000001110" when "011011000",
      "01101100110010110111001100100001001011000011010101000001010010101110000100000011010011000011110" when "011011001",
      "01101101010010111000111001000110111011001111011000000101000101110111011000100010100010001001010" when "011011010",
      "01101101110010111010100110001100101110110101001100011110110111001101111100111001110101101111100" when "011011011",
      "01101110010010111100010011110010100101110101110010011000110101110111011110101110011011011000000" when "011011100",
      "01101110110010111110000001111000100000010010001001111101010011111010010100101000111110110101010" when "011011101",
      "01101111010010111111110000011110011110001011010011010110100110011101011110100001101101010111111" when "011011110",
      "01101111110011000001011111100100011111100010001110101111000101101000100101101100011000111101110" when "011011111",
      "01110000010011000011001111001010100100010111111100010001001100100011111101000100011011100010000" when "011100000",
      "01110000110011000100111111010000101100101101011100000111011001011000100001011000111010001101011" when "011100001",
      "01110001010011000110101111110110111000100011101110011100001101001111111001011000101000100111110" when "011100010",
      "01110001110011001000100000111101000111111011110011011010001100010100010101111110001100001010110" when "011100011",
      "01110010010011001010010010100011011010110110101011001011111101110000110010011011111111010101110" when "011100100",
      "01110010110011001100000100101001110001010101010101111100001011110000110100101000010101000001001" when "011100101",
      "01110011010011001101110111010000001011011000110011110101100011100000101101001001011011110100110" when "011100110",
      "01110011110011001111101010010110101001000010000101000010110101001101010111100001100001011110001" when "011100111",
      "01110100010011010001011101111101001010010010001001101110110100000100011010011010110110000110110" when "011101000",
      "01110100110011010011010010000011101111001010000010000100010110010100000111110011101111101101011" when "011101001",
      "01110101010011010101000110101010010111101010101110001110010101001011011101001010101101011110101" when "011101010",
      "01110101110011010110111011110001000011110101001110010111101100111010000011101010011011001111001" when "011101011",
      "01110110010011011000110001010111110011101010100010101011011100110000010000010101110100110110110" when "011101100",
      "01110110110011011010100111011110100111001011101011010100100110111111000100010100001001101100000" when "011101101",
      "01110111010011011100011110000101011110011001101000011110010000111000001100111101000000000001100" when "011101110",
      "01110111110011011110010101001100011001010101011010010011100010101110000100000100011000100100000" when "011101111",
      "01111000010011100000001100110011011000000000000000111111100111110011110000000110110001111000100" when "011110000",
      "01111000110011100010000100111010011010011010011100101101101110011101000100010101001011111100001" when "011110001",
      "01111001010011100011111101100001100000100101101101101001000111111110100001000001001011100101010" when "011110010",
      "01111001110011100101110110101000101010100010110011111101001000101101010011101000111110000101000" when "011110011",
      "01111010010011100111110000001111111000010010101111110101000111111111010111000011011100101001001" when "011110100",
      "01111010110011101001101010010111001001110110100001011100100000001011010011101100010000000000101" when "011110101",
      "01111011010011101011100100111110011111001111001000111110101110101000011111101111110011111111010" when "011110110",
      "01111011110011101101100000000101111000011101100110100111010011101110111111010111011011000011100" when "011110111",
      "01111100010011101111011011101101010101100010111010100001110010110111100100110101010001111100100" when "011111000",
      "01111100110011110001010111110100110110100000000100111001110010011011110000110000100011010001100" when "011111001",
      "01111101010011110011010100011100011011010110000101111010111011110101110010010001011011001010010" when "011111010",
      "01111101110011110101010001100100000100000101111101110000111011100000100111001101001010111000000" when "011111011",
      "01111110010011110111001111001011110000110000101100100111100000110111111100010010001100011111100" when "011111100",
      "01111110110011111001001101010011100001010111010010101010011110011000001101010100000110100100000" when "011111101",
      "01111111010011111011001011111011010101111010110000000101101001011110100101010111101111110011101" when "011111110",
      "01111111110011111101001011000011001110011100000101000100111010101000111110111111010010110100000" when "011111111",
      "10000000000011111110001010110011001100001100010000011101110011111101101111101100101100001000100" when "100000000",
      "10000000100100000000001010101011001010101100010001001001100110101011111001101011111100001111101" when "100000001",
      "10000001000100000010001011000011001101001100101001110111011001110100001000011011110111111100001" when "100000010",
      "10000001100100000100001011111011010011101110011010110011010000010110111110000100001100101101011" when "100000011",
      "10000010000100000110001101010011011110010010100100001001010000010101101101000000001100110000100" when "100000100",
      "10000010100100001000001111001011101100111010000110000101100010110010011000001010110010110010000" when "100000101",
      "10000011000100001010010001100011111111100110000000110100010011101111110011001010100101110001000" when "100000110",
      "10000011100100001100010100011100010110010111010100100001110010010001100010011101111100110011011" when "100000111",
      "10000100000100001110010111110100110001001111000001011010010000011011111011100111000010111010100" when "100001000",
      "10000100100100010000011011101101010000001110000111101010000011010100000101010111111010111001001" when "100001001",
      "10000101000100010010100000000101110011010101100111011101100010111111110111111110100011001010011" when "100001010",
      "10000101100100010100100100111110011010100110100001000001001010100101111101010000111001101001100" when "100001011",
      "10000110000100010110101010010111000110000001110100100001011000001101110000111000111111101010101" when "100001100",
      "10000110100100011000110000001111110101101000100010001010101100111111100000100000111101110100000" when "100001101",
      "10000111000100011010110110101000101001011011101010001001101101000100001011111111000111111001010" when "100001110",
      "10000111100100011100111101100001100001011100001100101010111111100101100101100010000000110110100" when "100001111",
      "10001000000100011111000100111010011101101011001001111011001110101110010001111100011110101101001" when "100010000",
      "10001000100100100001001100110011011110001001100010000111000111101001101000110001101110100000110" when "100010001",
      "10001001000100100011010101001100100010111000010101011011011010100011110100100001011000010110011" when "100010010",
      "10001001100100100101011110000101101011111000100100000100111010101001110010110011100011010010110" when "100010011",
      "10001010000100100111100111011110111001001011001110010000011110001001010100100100111001011011100" when "100010100",
      "10001010100100101001110001011000001010110001010100001010111110010000111110010010101011110111111" when "100010101",
      "10001011000100101011111011110001100000101011110110000001010111010000001000000110110110110011001" when "100010110",
      "10001011100100101110000110101010111010111011110100000000101000010110111110000100000101011111010" when "100010111",
      "10001100000100110000010010000100011001100010001110010101110011110110100000010001110110011001100" when "100011000",
      "10001100100100110010011101111101111100100000000101001101111111000000100011001000011111001111000" when "100011001",
      "10001101000100110100101010010111100011110110011000110110010010000111101111011101010001000010111" when "100011010",
      "10001101100100110110110111010001001111100110001001011011111000011111100010101110011100010101000" when "100011011",
      "10001110000100111001000100101010111111110000010111001100000000011100001111001111010101001010001" when "100011100",
      "10001110100100111011010010100100110100010110000010010011111011010010111100010100010111010011111" when "100011101",
      "10001111000100111101100000111110101101011000001011000000111101011001100110011111001010011011100" when "100011110",
      "10001111100100111111101111111000101010110111110001100000011110000110111111101010100110001011110" when "100011111",
      "10010000000101000001111111010010101100110101110101111111110111110010101111010110110110011100100" when "100100000",
      "10010000100101000100001111001100110011010011011000101100100111110101010010110101011111011111111" when "100100001",
      "10010001000101000110011111100110111110010001011001110100001110100111111101010101100010001111001" when "100100010",
      "10010001100101001000110000100001001101110000111001100100001111100100111000001111100000011001001" when "100100011",
      "10010010000101001011000001111011100001110010111000001010010001000111000011010001100000110010001" when "100100100",
      "10010010100101001101010011110101111010011000010101110011111100101010010100101011010011100011100" when "100100101",
      "10010011000101001111100110010000010111100010010010101110111110101011011001011010010110011101110" when "100100110",
      "10010011100101010001111001001010111001010001101111001001000110100111110101010101111001001001110" when "100100111",
      "10010100000101010100001100100101011111100111101011010000000110111110000011011011000001011100110" when "100101000",
      "10010100100101010110100000100000001010100101000111010001110101001101010101111000101111101011111" when "100101001",
      "10010101000101011000110100111010111010001011000011011100001001110101110110011100000011000001011" when "100101010",
      "10010101100101011011001001110101101110011010011111111101000000011000100110011011111101110010110" when "100101011",
      "10010110000101011101011111010000100111010100011101000010010111010111011111000101101001110111011" when "100101100",
      "10010110100101011111110101001011100100111001111010111010010000010101010001101000011101000000100" when "100101101",
      "10010111000101100010001011100110100111001011111001110010101111110101100111100001111101010010001" when "100101110",
      "10010111100101100100100010100001101110001011011001111001111101011101000010101010000101011100100" when "100101111",
      "10011000000101100110111001111100111001111001011011011110000011110000111101011111001001010111001" when "100110000",
      "10011000100101101001010001111000001010010110111110101101010000010111101011010001111010011100010" when "100110001",
      "10011001000101101011101010010011011111100101000011110101110011111000011000010001101100000101001" when "100110010",
      "10011001100101101110000011001110111001100100101011000110000001111011001001111000011000001000011" when "100110011",
      "10011010000101110000011100101010011000010110110100101100010001001000111110110110100011010111100" when "100110100",
      "10011010100101110010110110100101111011111100100000110110111011001011101111011111100001111110111" when "100110101",
      "10011011000101110101010001000001100100010110101111110100011100101110001101110101011100000101110" when "100110110",
      "10011011100101110111101011111101010001100110100001110011010101011100000101110101010010010000001" when "100110111",
      "10011100000101111010000111011001000011101100110111000010001000000001111101100011000010000000010" when "100111000",
      "10011100100101111100100011010100111010101010101111101111011010001101010101010101101010011010011" when "100111001",
      "10011101000101111110111111110000110110100001001100001001110100101100101000000011010000101000100" when "100111010",
      "10011101100110000001011100101100110111010001001100100000000011001111001011001101000100011111111" when "100111011",
      "10011110000110000011111010001000111100111011110001000000110100100101001111001011100101000110011" when "100111100",
      "10011110100110000110011000000101000111100001111001111010111010011111111111011010100101011010011" when "100111101",
      "10011111000110001000110110100001010111000100100111011101001001110001100010100101010000111001110" when "100111110",
      "10011111100110001011010101011101101011100100111001110110011010001100111010110010010000001011001" when "100111111",
      "10100000000110001101110100111010000101000011110001010101100110100110000101101111101101101000000" when "101000000",
      "10100000100110010000010100110110100011100010001110001001101100110001111100111111011010000110110" when "101000001",
      "10100001000110010010110101010011000111000001010000100001101101100110010110000010110001100111001" when "101000010",
      "10100001100110010101010110001111101111100001111000101100101100111010000010100110111111111101111" when "101000011",
      "10100010000110010111110111101100011101000101000110111001110001100100110000110001000101100011101" when "101000100",
      "10100010100110011010011001101001001111101011111011011000000101011111001011001001111100000010010" when "101000101",
      "10100011000110011100111100000110000111010111010110010110110101100010111001001010011011000100111" when "101000110",
      "10100011100110011111011111000011000100001000011000000101010001101010011111000111011101001000010" when "101000111",
      "10100100000110100010000010100000000110000000000000110010101100110001011110011110000100001011110" when "101001000",
      "10100100100110100100100110011101001100111111010000101110011100110100010101111111011110100100011" when "101001001",
      "10100101000110100111001010111010011001000111001000000111111010110000100001111101001011101111011" when "101001010",
      "10100101100110101001101111110111101010011000100111001110100010100100011100010101000001000110101" when "101001011",
      "10100110000110101100010101010101000000110100101110010001110011001111011100111101001110110101110" when "101001100",
      "10100110100110101110111011010010011100011100011101100001001110110001111001110000100100110000001" when "101001101",
      "10100111000110110001100001101111111101010000110101001100011010001101000110111010010111001000010" when "101001110",
      "10100111100110110100001000101101100011010010110101100010111101100011010111000010100011100111010" when "101001111",
      "10101000000110110110110000001011001110100011011110110100100011110111111011011001110110000110000" when "101010000",
      "10101000100110111001011000001000111111000011110001010000111011001111000100000101101101100110111" when "101010001",
      "10101001000110111100000000100110110100110100101101000111110100101110000000001100100001010000111" when "101010010",
      "10101001100110111110101001100100101111110111010010101001000100011010111110000001100101001010111" when "101010011",
      "10101010000111000001010011000010110000001100100010000100100001011101001011010001001111011000101" when "101010100",
      "10101010100111000011111101000000110101110101011011101010000101111100110101001100111100111000100" when "101010101",
      "10101011000111000110100111011111000000110010111111101001101111000011001000110111010110100001100" when "101010110",
      "10101011100111001001010010011101010001000110001110010011011100111010010011010000010110000011101" when "101010111",
      "10101100000111001011111101111011100110110000000111110111010010101101100001100001001011000111100" when "101011000",
      "10101100100111001110101001111010000001110001101100100101010110101001000001001000100000010000011" when "101011001",
      "10101101000111010001010110011000100010001011111100101101110001111010000000000110011111111110010" when "101011010",
      "10101101100111010100000011010111000111111111111000100000110000101110101101001000111001110001010" when "101011011",
      "10101110000111010110110000110101110011001110100000001110100010010110010111110111000111001101100" when "101011100",
      "10101110100111011001011110110100100011111000110100000111011001000001010000111110010001000001000" when "101011101",
      "10101111000111011100001101010011011001111111110100011011101010000000101010011101010100001001011" when "101011110",
      "10101111100111011110111100010010010101100100100001011011101101100110110111110001000110111010110" when "101011111",
      "10110000000111100001101011110001010110100111111011010111111111000111001110000000011110001000010" when "101100000",
      "10110000100111100100011011110000011101001011000010100000111100110110000100001000010010001100011" when "101100001",
      "10110001000111100111001100001111101001001110110111000111001000001000110011000111100100010011110" when "101100010",
      "10110001100111101001111101001110111010110100011001011011000101010101110110001011100011100111001" when "101100011",
      "10110010000111101100101110101110010001111100101001101101011011110100101010111011110010010111101" when "101100100",
      "10110010100111101111100000101101101110101000101000001110110101111101110001100110001011001011101" when "101100101",
      "10110011000111110010010011001101010000111001010101010000000001001010101101001011000110001100000" when "101100110",
      "10110011100111110101000110001100111000101111110001000001101101110110000011101001011110010011010" when "101100111",
      "10110100000111110111111001101100100110001100111011110100101111011011011110001010110110011100101" when "101101000",
      "10110100100111111010101101101100011001010001110101111001111100010111101001001111011110110101001" when "101101001",
      "10110101000111111101100010001100010001111111011111100010001110001000010100111010011010001100100" when "101101010",
      "10110101101000000000010111001100010000010110111000111110100001001100010100111101100011001000001" when "101101011",
      "10110110001000000011001100101100010100011001000010011111110101000011100001000101110001010110001" when "101101100",
      "10110110101000000110000010101100011110000110111100010111001100001110110101000110111111000001101" when "101101101",
      "10110111001000001000111001001100101101100001100110110101101100010000010001001000001110001000000" when "101101110",
      "10110111101000001011110000001101000010101010000010001100011101101010111001101111101101101111100" when "101101111",
      "10111000001000001110100111101101011101100001001110101100101100000010111000001110111111011110000" when "101110000",
      "10111000101000010001011111101101111110001000001100100111100101111101011010101110111100110000110" when "101110001",
      "10111001001000010100011000001110100100011111111100001110011101000000110100011011111100010110100" when "101110010",
      "10111001101000010111010001001111010000101001011101110010100101110100011101110001110111101000011" when "101110011",
      "10111010001000011010001010110000000010100101110001100101011000000000110100101000010000000101011" when "101110100",
      "10111010101000011101000100110000111010010101110111111000001110001111011100011110010100101110000" when "101110101",
      "10111011001000011111111111010001110111111010110000111100100110001010111110100111000111100001101" when "101110110",
      "10111011101000100010111010010010111011010101011101000100000000011111001010010101100010111011010" when "101110111",
      "10111100001000100101110101110100000100100110111100100000000000111000110101001000011111010001010" when "101111000",
      "10111100101000101000110001110101010011110000001111100010001110000101111010110110111000010100100" when "101111001",
      "10111101001000101011101110010110101000110010010110011100010001110101011101111011110010110000111" when "101111010",
      "10111101101000101110101011011000000011101110010001011111111000110111100111100010100001101111010" when "101111011",
      "10111110001000110001101000111001100100100101000000111110110010111101100111110010101100010111101" when "101111100",
      "10111110101000110100100110111011001011010111100101001010110010111001110101111100010011010100100" when "101111101",
      "10111111001000110111100101011100111000000110111110010101101110011111110000100011110110010111110" when "101111110",
      "10111111101000111010100100011110101010110100001100110001011110100011111101101110011001111111100" when "101111111",
      "11000000001000111101100100000000100011100000010000101111111110111100001011001101101100111100100" when "110000000",
      "11000000101001000000100100000010100010001100001010100011001110011111001110101100001101111001011" when "110000001",
      "11000001001001000011100100100100100110111000111010011101001111000101000101111001010001000011000" when "110000010",
      "11000001101001000110100101100110110001100111100000110000000101100110110110110101000101110001010" when "110000011",
      "11000010001001001001100111001001000010011000111101101101111001111110101111111100111100010001010" when "110000100",
      "11000010101001001100101001001011011001001110010001101000110111001000001000010111001011010000100" when "110000101",
      "11000011001001001111101011101101110110001000011100110011001010111111011111111111010101101000101" when "110000110",
      "11000011101001010010101110110000011001001000011111011111000110100010011111110010010000001100010" when "110000111",
      "11000100001001010101110010010011000010001111011001111110111101101111111001111010000111010101000" when "110001000",
      "11000100101001011000110110010101110001011110001100100101000111100111101001111010100100110010011" when "110001001",
      "11000101001001011011111010111000100110110101110111100011111110001010110100111100110101011001001" when "110001010",
      "11000101101001011110111111111011100010010111011011001101111110011011101001111011101110110100001" when "110001011",
      "11000110001001100010000101011110100100000011110111110101101000011101100001101111110101010110010" when "110001100",
      "11000110101001100101001011100001101011111100001101101101011111010100111111011011100001101100101" when "110001101",
      "11000111001001101000010010000100111010000001011101001000001001000111110000010111000110110010001" when "110001110",
      "11000111101001101011011001001000001110010100100110011000001110111100101100011100110111100100001" when "110001111",
      "11001000001001101110100000101011101000110110101001110000011100111011110110010101001100110111100" when "110010000",
      "11001000101001110001101000101111001001101000100111100011100010001110011011100010101011001111100" when "110010001",
      "11001001001001110100110001010010110000101011100000000100010000111110110100101110001000110100110" when "110010010",
      "11001001101001110111111010010110011110000000010011100101011110011000100101110010110011001101010" when "110010011",
      "11001010001001111011000011111010010001101000000010011010000010101000011110001010010101010110001" when "110010100",
      "11001010101001111110001101111110001011100011101100110100111000111100011000111000111101011101010" when "110010101",
      "11001011001010000001011000100010001011110100010011001000111111100011011100111001100010111101000" when "110010110",
      "11001011101010000100100011100110010010011010110101101001010111101101111101001001101100010111011" when "110010111",
      "11001100001010000111101111001010011111011000010100101001000101101101011000110101110101010011110" when "110011000",
      "11001100101010001010111011001110110010101101110000011011010000110100011011100101010100011100100" when "110011001",
      "11001101001010001110000111110011001100011100001001010011000011010110111101100110100001011101110" when "110011010",
      "11001101101010010001010100110111101100100100011111100011101010101010000011111010111011000101100" when "110011011",
      "11001110001010010100100010011100010011000111110011100000010111000100000000100011001101000100001" when "110011100",
      "11001110101010010111110000100001000000000111000101011100011011111100010010101011010110001110001" when "110011101",
      "11001111001010011010111111000101110011100011010101101011001111101011100110110110101110011111010" when "110011110",
      "11001111101010011110001110001010101101011101100100100000001011101011110111001100001100111101000" when "110011111",
      "11010000001010100001011101101111101101110110110010001110101100011000001011100010001101111100101" when "110100000",
      "11010000101010100100101101110100110100101111111111001010010001001100111001101010111001000111010" when "110100001",
      "11010001001010100111111110011010000010001010001011100110011100100111100101100000000111100001100" when "110100010",
      "11010001101010101011001111011111010110000110010111110110110100000111000001001111101001110001111" when "110100011",
      "11010010001010101110100001000100110000100101100100001111000000001011001101100111001110001001110" when "110100100",
      "11010010101010110001110011001010010001101000110001000010101100010101011010000000100110101110011" when "110100101",
      "11010011001010110101000101101111111001010000111110100101100111001000000100101101101111100011100" when "110100110",
      "11010011101010111000011000110101100111011111001101001011100010000110111011000100110100110101110" when "110100111",
      "11010100001010111011101100011011011100010100011101001000010001110110111001101100011001000111100" when "110101000",
      "11010100101010111111000000100001010111110001101110101111101101111110001100100111011011011101110" when "110101001",
      "11010101001011000010010101000111011001111000000010010101110001000100001111100001011101101101111" when "110101010",
      "11010101101011000101101010001101100010101000011000001110011000110001101101111010101010101100111" when "110101011",
      "11010110001011001000111111110011110010000011110000101101100101110000100011010011111100011111010" when "110101100",
      "11010110101011001100010101111010001000001011001100000111011011101011111011011011000010101001110" when "110101101",
      "11010111001011001111101100100000100100111111101010110000000001010000010010010110101000100011010" when "110101110",
      "11010111101011010011000011100111001000100010001100111011100000001011010100110010011011100111010" when "110101111",
      "11011000001011010110011011001101110010110011110010111110000101001100000000001011010001101010010" when "110110000",
      "11011000101011011001110011010100100011110101011101001100000000000010100010111011001111001101101" when "110110001",
      "11011001001011011101001011111011011011101000001011111001100011100000011100100101101101110101100" when "110110010",
      "11011001101011100000100101000010011010001100111111011011000101011000011110000011100010011111011" when "110110011",
      "11011010001011100011111110101001011111100100111000000100111110011110101001101111000011111001110" when "110110100",
      "11011010101011100111011000110000101011110000110110001011101010101000010011110000010000111100001" when "110110101",
      "11011011001011101010110011010111111110110001111010000011101000101100000010001000110111000000100" when "110110110",
      "11011011101011101110001110011111011000101001000100000001011010100001101101000000011000011110010" when "110110111",
      "11011100001011110001101010000110111001010111010100011001100101000010011110110000010011000100100" when "110111000",
      "11011100101011110101000110001110100000111101101011100000110000001000110100010000000110010111000" when "110111001",
      "11011101001011111000100010110110001111011101001001101011100110110000011101000001011010001011001" when "110111010",
      "11011101101011111011111111111110000100110110101111001110110110110110011011011100000101000101110" when "110111011",
      "11011110001011111111011101100110000001001011011100011111010001011001000100111010010010111010110" when "110111100",
      "11011110101100000010111011101110000100011100010001110001101010011000000010000100101011001100110" when "110111101",
      "11011111001100000110011010010110001110101010001111011010111000110100001110111110010111101101110" when "110111110",
      "11011111101100001001111001011110011111110110010101101111110110101111111011010001001011000001101" when "110111111",
      "11100000001100001101011001000110111000000001100101000101100001001110101010011001100111000000111" when "111000000",
      "11100000101100010000111001001111010111001100111101110000111000010101010011110011000011011011111" when "111000001",
      "11100001001100010100011001110111111101011001100000000110111111001010000011000011110100100000011" when "111000010",
      "11100001101100010111111011000000101010101000001100011100111011110100011000001001010001011110100" when "111000011",
      "11100010001100011011011100101001011110111010000011000111110111011101000111100011111011001111111" when "111000100",
      "11100010101100011110111110110010011010010000000100011100111110001110011010100011100010111110111" when "111000101",
      "11100011001100100010100001011011011100101011010000110001011111010011101111010011010000101111100" when "111000110",
      "11100011101100100110000100100100100110001100101000011010101100111001111001000101101010001000100" when "111000111",
      "11100100001100101001101000001101110110110101001011101101111100001111000000100000111000111110000" when "111001000",
      "11100100101100101101001100010111001110100101111011000000100101100010100011101010110001111101000" when "111001001",
      "11100101001100110000110001000000101101011111110110101000000100000101010110010100111011010111010" when "111001010",
      "11100101101100110100010110001010010011100011111110111001110110001001100010001000110011110001000" when "111001011",
      "11100110001100110111111011110100000000110011010100001011011101000010100110110011111000101110111" when "111001100",
      "11100110101100111011100001111101110101001110110110110010011101000101011010010011101101100101010" when "111001101",
      "11100111001100111111001000100111110000110111100111000100011101101000001001000010000010001000010" when "111001110",
      "11100111101101000010101111110001110011101110100101010111001001000010010110000000111001011100110" when "111001111",
      "11101000001101000110010111011011111101110100110010000000001100101100111011000110110000101010101" when "111010000",
      "11101000101101001001111111100110001111001011001101010101011001000010001001001010100101101111011" when "111010001",
      "11101001001101001101101000010000100111110010110111101100100001011101101000001111111110010010010" when "111010010",
      "11101001101101010001010001011011000111101100110001011011011100011100010111110011001110011001001" when "111010011",
      "11101010001101010100111011000101101110111001111010111000000011011100101110110101011111011101111" when "111010100",
      "11101010101101011000100101010000011101011011010100011000010010111110011100001000110111000110000" when "111010101",
      "11101011001101011100001111111011010011010001111110010010001010100010100110011100011101111001001" when "111010110",
      "11101011101101011111111011000110010000011110111000111011101100101011101100101000100110011010101" when "111010111",
      "11101100001101100011100110110001010101000011000100101010111110111101100101111010110100000010111" when "111011000",
      "11101100101101100111010010111100100000111111100001110110001001111101100010000010000001111001100" when "111011001",
      "11101101001101101010111111100111110100010101010000110011011001010010001001011010101001110001011" when "111011010",
      "11101101101101101110101100110011001111000101010001111000111011100011011101011010101011000100101" when "111011011",
      "11101110001101110010011010011110110001010000100101011101000010011010111000011101110001110010001" when "111011100",
      "11101110101101110110001000101010011010111000001011110110000010100011001110010001011101011011111" when "111011101",
      "11101111001101111001110111010110001011111101000101011010010011101000101100000001001000000110100" when "111011110",
      "11101111101101111101100110100010000100100000010010100000010000011000111000100010001101011000111" when "111011111",
      "11110000001110000001010110001110000100100010110011011110010110100010110100100000010001011101101" when "111100000",
      "11110000101110000101000110011010001100000101101000101011000110110110111010101001001000000101101" when "111100001",
      "11110001001110001000110111000110011011001001110010011101000101000110111111111000111011101010001" when "111100010",
      "11110001101110001100101000010010110001110000010001001010111000000110010011100110010100010010000" when "111100011",
      "11110010001110010000011001111111001111111010000101001011001001101001011111101110011110110101010" when "111100100",
      "11110010101110010100001100001011110101101000001110110100100110100110101001000001010100000100011" when "111100101",
      "11110011001110010111111110111000100010111011101110011101111110110101001111001101011111101110000" when "111100110",
      "11110011101110011011110010000101010111110101100100011110000101001110001101001100100111100111100" when "111100111",
      "11110100001110011111100101110010010100010110110001001011101111101011111001001111010010110101010" when "111101000",
      "11110100101110100011011001111111011000100000010100111101110111001010000101001001010000110100110" when "111101001",
      "11110101001110100111001110101100100100010011010000001011010111100101111110011101100000100110110" when "111101010",
      "11110101101110101011000011111001110111110000100011001011001111111110001110101010010111111011100" when "111101011",
      "11110110001110101110111001100111010010111001001110010100100010010010111011010101101010011110101" when "111101100",
      "11110110101110110010101111110100110101101110010001111110010011100101100110011000110001000100111" when "111101101",
      "11110111001110110110100110100010100000010000101110011111101011111001001110001100110000111010111" when "111101110",
      "11110111101110111010011101110000010010100001100100001111110110010010001101110110100010110100001" when "111101111",
      "11111000001110111110010101011110001100100001110011100110000000110110011101010010111010011011001" when "111110000",
      "11111000101111000010001101101100001110010010011100111001011100101101010001100010101101100011100" when "111110001",
      "11111001001111000110000110011010010111110100100000100001011101111111011100110110111011011011010" when "111110010",
      "11111001101111001001111111101000101001001000111110110101011011110111001110111100110011111110101" when "111110011",
      "11111010001111001101111001010111000010010000111000001100110000100000010101001001111111001011111" when "111110100",
      "11111010101111010001110011100101100011001101001100111110111001000111111010101000100100011000100" when "111110101",
      "11111011001111010101101110010100001011111110111101100011010101111100101000100011010001100111010" when "111110110",
      "11111011101111011001101001100010111100100111001010010001101010001110100110010001100010111111000" when "111110111",
      "11111100001111011101100101010001110101000110110011100001011100001111011001100011101010000010111" when "111111000",
      "11111100101111100001100001100000110101011110111001101010010101010010000110101110110101001010110" when "111111001",
      "11111101001111100101011110001111111101110000011101000100000001101011010000111001010110111101011" when "111111010",
      "11111101101111101001011011011111001101111100011110000110010000110000111010000110101101101011001" when "111111011",
      "11111110001111101101011001001110100110000011111101001000110100111010100011100011101010101001101" when "111111100",
      "11111110101111110001010111011110000110000111111010100011100011100001001101110010011001110000011" when "111111101",
      "11111111001111110101010110001101101110001001010110101110010100111111011000110110101000110110011" when "111111110",
      "11111111101111111001010101011101011110001001010010000001000100110001000100100001101111010000111" when "111111111",
      "-----------------------------------------------------------------------------------------------" when others;
   Y1_c2 <= Y0_c2; -- for the possible blockram register
   Y <= Y1_c2;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_104_Freq300_uid43
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_104_Freq300_uid43 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(103 downto 0);
          Y : in  std_logic_vector(103 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(103 downto 0)   );
end entity;

architecture arch of IntAdder_104_Freq300_uid43 is
signal Rtmp_c2 :  std_logic_vector(103 downto 0);
signal X_c1, X_c2 :  std_logic_vector(103 downto 0);
signal Cin_c1, Cin_c2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               X_c1 <= X;
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               X_c2 <= X_c1;
               Cin_c2 <= Cin_c1;
            end if;
         end if;
      end process;
   Rtmp_c2 <= X_c2 + Y + Cin_c2;
   R <= Rtmp_c2;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable2_Freq300_uid45
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable2_Freq300_uid45 is
    port (clk, ce_4 : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(86 downto 0)   );
end entity;

architecture arch of LogTable2_Freq300_uid45 is
signal Y0_c4 :  std_logic_vector(86 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c4 :  std_logic_vector(86 downto 0);
signal X_c4 :  std_logic_vector(8 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_4 = '1' then
               X_c4 <= X;
            end if;
         end if;
      end process;
   with X_c4  select  Y0_c4 <= 
      "000000000000000000000000000000000000000000000000000011111111111111111111111111111111111" when "000000000",
      "000000001000000000000000000000000000111111100000000100000000001010100010101100101010100" when "000000001",
      "000000010000000000000000000000000011111111000000000100000001010100110101011001010101101" when "000000010",
      "000000011000000000000000000000001000111110100000000100000100011110111000000110000010011" when "000000011",
      "000000100000000000000000000000001111111110000000000100001010101000101010110010110010100" when "000000100",
      "000000101000000000000000000000011000111101100000000100010100110010001101011111101000101" when "000000101",
      "000000110000000000000000000000100011111101000000000100100011111011100000001100101000010" when "000000110",
      "000000111000000000000000000000110000111100100000000100111001000100100010111001110101011" when "000000111",
      "000001000000000000000000000000111111111100000000000101010101001101010101100111010100111" when "000001000",
      "000001001000000000000000000001010000111011100000000101111001010101111000010101001100100" when "000001001",
      "000001010000000000000000000001100011111011000000000110100110011110001011000011100010100" when "000001010",
      "000001011000000000000000000001111000111010100000000111011101100110001101110010011110000" when "000001011",
      "000001100000000000000000000010001111111010000000001000011111101110000000100010000111000" when "000001100",
      "000001101000000000000000000010101000111001100000001001101101110101100011010010100110000" when "000001101",
      "000001110000000000000000000011000011111001000000001011001000111100110110000100000100011" when "000001110",
      "000001111000000000000000000011100000111000100000001100110010000011111000110110101100010" when "000001111",
      "000010000000000000000000000011111111111000000000001110101010001010101011101010101000100" when "000010000",
      "000010001000000000000000000100100000110111100000010000110010010001001110100000000100110" when "000010001",
      "000010010000000000000000000101000011110111000000010011001011010111100001010111001101100" when "000010010",
      "000010011000000000000000000101101000110110100000010101110110011101100100010000001111110" when "000010011",
      "000010100000000000000000000110001111110110000000011000110100100011010111001011011001010" when "000010100",
      "000010101000000000000000000110111000110101100000011100000110101000111010001000111000111" when "000010101",
      "000010110000000000000000000111100011110101000000011111101101101110001101001000111101110" when "000010110",
      "000010111000000000000000001000010000110100100000100011101010110011010000001011111000010" when "000010111",
      "000011000000000000000000001000111111110100000000100111111110111000000011010001111001001" when "000011000",
      "000011001000000000000000001001110000110011100000101100101010111100100110011011010001111" when "000011001",
      "000011010000000000000000001010100011110011000000110001110000000000111001101000010101001" when "000011010",
      "000011011000000000000000001011011000110010100000110111001111000100111100111001010101110" when "000011011",
      "000011100000000000000000001100001111110010000000111101001001001000110000001110100111110" when "000011100",
      "000011101000000000000000001101001000110001100001000011011111001100010011101000011111110" when "000011101",
      "000011110000000000000000001110000011110001000001001010010010001111100111000111010011001" when "000011110",
      "000011111000000000000000001111000000110000100001010001100011010010101010101011011000000" when "000011111",
      "000100000000000000000000001111111111110000000001011001010011010101011110010101000101010" when "000100000",
      "000100001000000000000000010001000000101111100001100001100011011000000010000100110010011" when "000100001",
      "000100010000000000000000010010000011101111000001101010010100011010010101111010110111111" when "000100010",
      "000100011000000000000000010011001000101110100001110011100111011100011001110111101110110" when "000100011",
      "000100100000000000000000010100001111101110000001111101011101011110001101111011110001001" when "000100100",
      "000100101000000000000000010101011000101101100010000111110111011111110010000111011001011" when "000100101",
      "000100110000000000000000010110100011101101000010010010110110100001000110011011000010111" when "000100110",
      "000100111000000000000000010111110000101100100010011110011011100010001010110111001010000" when "000100111",
      "000101000000000000000000011000111111101100000010101010100111100010111111011100001011010" when "000101000",
      "000101001000000000000000011010010000101011100010110111011011100011100100001010100100101" when "000101001",
      "000101010000000000000000011011100011101011000011000100111000100011111001000010110100010" when "000101010",
      "000101011000000000000000011100111000101010100011010010111111100011111110000101011001010" when "000101011",
      "000101100000000000000000011110001111101010000011100001110001100011110011010010110011101" when "000101100",
      "000101101000000000000000011111101000101001100011110001001111100011011000101011100100000" when "000101101",
      "000101110000000000000000100001000011101001000100000001011010100010101110010000001011100" when "000101110",
      "000101111000000000000000100010100000101000100100010010010011100001110100000001001100101" when "000101111",
      "000110000000000000000000100011111111101000000100100011111011100000101001111111001010000" when "000110000",
      "000110001000000000000000100101100000100111100100110110010011011111010000001010100111010" when "000110001",
      "000110010000000000000000100111000011100111000101001001011100011101100110100100001000110" when "000110010",
      "000110011000000000000000101000101000100110100101011101010111011011101101001100010011110" when "000110011",
      "000110100000000000000000101010001111100110000101110010000101011001100100000011101110000" when "000110100",
      "000110101000000000000000101011111000100101100110000111100111010111001011001010111110001" when "000110101",
      "000110110000000000000000101101100011100101000110011101111110010100100010100010101011101" when "000110110",
      "000110111000000000000000101111010000100100100110110101001011010001101010001011011110100" when "000110111",
      "000111000000000000000000110000111111100100000111001101001111001110100010000101111111101" when "000111000",
      "000111001000000000000000110010110000100011100111100110001011001011001010010010111000101" when "000111001",
      "000111010000000000000000110100100011100011001000000000000000000111100010110010110100000" when "000111010",
      "000111011000000000000000110110011000100010101000011010101111000011101011100110011100110" when "000111011",
      "000111100000000000000000111000001111100010001000110110011000111111100100101110011110101" when "000111100",
      "000111101000000000000000111010001000100001101001010010111110111011001110001011100110100" when "000111101",
      "000111110000000000000000111100000011100001001001110000100001110110100111111110100001101" when "000111110",
      "000111111000000000000000111110000000100000101010001111000010110001110010000111111110001" when "000111111",
      "001000000000000000000000111111111111100000001010101110100010101100101100101000101010111" when "001000000",
      "001000001000000000000001000010000000011111101011001111000010100111010111100001010111100" when "001000001",
      "001000010000000000000001000100000011011111001011110000100011100001110010110010110100100" when "001000010",
      "001000011000000000000001000110001000011110101100010011000110011011111110011101110010110" when "001000011",
      "001000100000000000000001001000001111011110001100110110101100010101111010100011000100010" when "001000100",
      "001000101000000000000001001010011000011101101101011011010110001111100111000011011011100" when "001000101",
      "001000110000000000000001001100100011011101001110000001000101001001000011111111101100001" when "001000110",
      "001000111000000000000001001110110000011100101110100111111010000010010001011000101010001" when "001000111",
      "001001000000000000000001010000111111011100001111001111110101111011001111001111001010010" when "001001000",
      "001001001000000000000001010011010000011011101111111000111001110011111101100100000010011" when "001001001",
      "001001010000000000000001010101100011011011010000100011000110101100011100011000001000101" when "001001010",
      "001001011000000000000001010111111000011010110001001110011101100100101011101100010100010" when "001001011",
      "001001100000000000000001011010001111011010010001111010111111011100101011100001011101001" when "001001100",
      "001001101000000000000001011100101000011001110010101000101101010100011011111000011011110" when "001001101",
      "001001110000000000000001011111000011011001010011010111101000001011111100110010001001110" when "001001110",
      "001001111000000000000001100001100000011000110100000111110001000011001110001111100001000" when "001001111",
      "001010000000000000000001100011111111011000010100111001001000111010010000010001011100011" when "001010000",
      "001010001000000000000001100110100000010111110101101011110000110001000010111000110111110" when "001010001",
      "001010010000000000000001101001000011010111010110011111101001100111100110000110101111010" when "001010010",
      "001010011000000000000001101011101000010110110111010100110100011101111001111100000000000" when "001010011",
      "001010100000000000000001101110001111010110011000001011010010010011111110011001101000000" when "001010100",
      "001010101000000000000001110000111000010101111001000011000100001001110011100000100101111" when "001010101",
      "001010110000000000000001110011100011010101011001111100001010111111011001010001111000111" when "001010110",
      "001010111000000000000001110110010000010100111010110110100111110100101111101110100001010" when "001010111",
      "001011000000000000000001111000111111010100011011110010011011101001110110110111011111110" when "001011000",
      "001011001000000000000001111011110000010011111100101111100111011110101110101101110110000" when "001011001",
      "001011010000000000000001111110100011010011011101101110001100010011010111010010100110101" when "001011010",
      "001011011000000000000010000001011000010010111110101110001011000111110000100110110100100" when "001011011",
      "001011100000000000000010000100001111010010011111101111100100111011111010101011100011100" when "001011100",
      "001011101000000000000010000111001000010010000000110010011010101111110101100001111000010" when "001011101",
      "001011110000000000000010001010000011010001100001110110101101100011100001001010111000010" when "001011110",
      "001011111000000000000010001101000000010001000010111100011110010110111101100111101001100" when "001011111",
      "001100000000000000000010001111111111010000100100000011101110001010001010111001010010111" when "001100000",
      "001100001000000000000010010011000000010000000101001100011101111101001001000000111100001" when "001100001",
      "001100010000000000000010010110000011001111100110010110101110101111110111111111101101100" when "001100010",
      "001100011000000000000010011001001000001111000111100010100001100010010111110110110000001" when "001100011",
      "001100100000000000000010011100001111001110101000101111110111010100101000100111001110000" when "001100100",
      "001100101000000000000010011111011000001110001001111110110001000110101010010010010001100" when "001100101",
      "001100110000000000000010100010100011001101101011001111001111111000011100111001000110010" when "001100110",
      "001100111000000000000010100101110000001101001100100001010100101010000000011100111000010" when "001100111",
      "001101000000000000000010101000111111001100101101110101000000011011010100111110110100100" when "001101000",
      "001101001000000000000010101100010000001100001111001010010100001100011010100000001000011" when "001101001",
      "001101010000000000000010101111100011001011110000100001010000111101010001000010000010100" when "001101010",
      "001101011000000000000010110010111000001011010001111001110111101101111000100101110001110" when "001101011",
      "001101100000000000000010110110001111001010110011010100001001011110010001001100100110010" when "001101100",
      "001101101000000000000010111001101000001010010100110000000111001110011010110111110000100" when "001101101",
      "001101110000000000000010111101000011001001110110001101110001111110010101101000100001110" when "001101110",
      "001101111000000000000011000000100000001001010111101101001010101110000001100000001100011" when "001101111",
      "001110000000000000000011000011111111001000111001001110010010011101011110100000000011001" when "001110000",
      "001110001000000000000011000111100000001000011010110001001010001100101100101001011001100" when "001110001",
      "001110010000000000000011001011000011000111111100010101110010111011101011111101100100001" when "001110010",
      "001110011000000000000011001110101000000111011101111100001101101010011100011101111000000" when "001110011",
      "001110100000000000000011010010001111000110111111100100011011011000111110001011101010111" when "001110100",
      "001110101000000000000011010101111000000110100001001110011101000111010001001000010011100" when "001110101",
      "001110110000000000000011011001100011000110000010111010010011110101010101010101001001010" when "001110110",
      "001110111000000000000011011101010000000101100100101000000000100011001010110011100100010" when "001110111",
      "001111000000000000000011100000111111000101000110010111100100010000110001100100111101011" when "001111000",
      "001111001000000000000011100100110000000100101000001000111111111110001001101010101110010" when "001111001",
      "001111010000000000000011101000100011000100001001111100010100101011010011000110010001001" when "001111010",
      "001111011000000000000011101100011000000011101011110001100011011000001101111001000001010" when "001111011",
      "001111100000000000000011110000001111000011001101101000101101000100111010000100011010100" when "001111100",
      "001111101000000000000011110100001000000010101111100001110010110001010111101001111001100" when "001111101",
      "001111110000000000000011111000000011000010010001011100110101011101100110101010111011100" when "001111110",
      "001111111000000000000011111100000000000001110011011001110110001001100111001000111110110" when "001111111",
      "010000000000000000000011111111111111000001010101011000110101110101011001000101100010000" when "010000000",
      "010000001000000000000100000100000000000000110111011001110101100000111100100010000101000" when "010000001",
      "010000010000000000000100001000000011000000011001011100110110001100010001100000001000001" when "010000010",
      "010000011000000000000100001100000111111111111011100001111000110111011000000001001100100" when "010000011",
      "010000100000000000000100010000001110111111011101101000111110100010010000000110110011110" when "010000100",
      "010000101000000000000100010100010111111110111111110010001000001100111001110010100000110" when "010000101",
      "010000110000000000000100011000100010111110100001111101010110110111010101000101110111000" when "010000110",
      "010000111000000000000100011100101111111110000100001010101011100001100010000010011010010" when "010000111",
      "010001000000000000000100100000111110111101100110011010000111001011100000101001101111101" when "010001000",
      "010001001000000000000100100101001111111101001000101011101010110101010000111101011100110" when "010001001",
      "010001010000000000000100101001100010111100101010111111010111011110110010111111000111110" when "010001010",
      "010001011000000000000100101101110111111100001101010101001110001000000110110000011000000" when "010001011",
      "010001100000000000000100110010001110111011101111101101001111110001001100010010110101100" when "010001100",
      "010001101000000000000100110110100111111011010010000111011101011010000011101000001000100" when "010001101",
      "010001110000000000000100111011000010111010110100100011111000000010101100110001111010100" when "010001110",
      "010001111000000000000100111111011111111010010111000010100000101011000111110001110101110" when "010001111",
      "010010000000000000000101000011111110111001111001100011011000010011010100101001100101000" when "010010000",
      "010010001000000000000101001000011111111001011100000110011111111011010011011010110011111" when "010010001",
      "010010010000000000000101001101000010111000111110101011111000100011000100000111001110110" when "010010010",
      "010010011000000000000101010001100111111000100001010011100011001010100110110000100011000" when "010010011",
      "010010100000000000000101010110001110111000000011111101100000110001111011011000011110001" when "010010100",
      "010010101000000000000101011010110111110111100110101001110010011001000010000000101111000" when "010010101",
      "010010110000000000000101011111100010110111001001011000011000111111111010101011000100110" when "010010110",
      "010010111000000000000101100100001111110110101100001001010101100110100101011001001111110" when "010010111",
      "010011000000000000000101101000111110110110001110111100101001001101000010001101000000110" when "010011000",
      "010011001000000000000101101101101111110101110001110010010100110011010001001000001001011" when "010011001",
      "010011010000000000000101110010100010110101010100101010011001011001010010001100011100000" when "010011010",
      "010011011000000000000101110111010111110100110111100100110111111111000101011011101011110" when "010011011",
      "010011100000000000000101111100001110110100011010100001110001100100101010110111101100101" when "010011100",
      "010011101000000000000110000001000111110011111101100001000111001010000010100010010011000" when "010011101",
      "010011110000000000000110000110000010110011100000100010111001101111001100011101010100100" when "010011110",
      "010011111000000000000110001010111111110011000011100111001010010100001000101010100111000" when "010011111",
      "010100000000000000000110001111111110110010100110101101111001111000110111001100000001101" when "010100000",
      "010100001000000000000110010100111111110010001001110111001001011101011000000011011011110" when "010100001",
      "010100010000000000000110011010000010110001101101000010111010000001101011010010101110000" when "010100010",
      "010100011000000000000110011111000111110001010000010001001100100101110000111011110001011" when "010100011",
      "010100100000000000000110100100001110110000110011100010000010001001101001000000011111101" when "010100100",
      "010100101000000000000110101001010111110000010110110101011011101101010011100010110011100" when "010100101",
      "010100110000000000000110101110100010101111111010001011011010010000110000100100101000100" when "010100110",
      "010100111000000000000110110011101111101111011101100011111110110100000000000111111010100" when "010100111",
      "010101000000000000000110111000111110101111000000111111001010010111000010001110100110100" when "010101000",
      "010101001000000000000110111110001111101110100100011100111101111001110110111010101010001" when "010101001",
      "010101010000000000000111000011100010101110000111111101011010011100011110001110000011110" when "010101010",
      "010101011000000000000111001000110111101101101011100000100000111110111000001010110010011" when "010101011",
      "010101100000000000000111001110001110101101001111000110010010100001000100110010110110000" when "010101100",
      "010101101000000000000111010011100111101100110010101110110000000011000100001000001111010" when "010101101",
      "010101110000000000000111011001000010101100010110011001111010100100110110001100111111100" when "010101110",
      "010101111000000000000111011110011111101011111010000111110011000110011011000011001000111" when "010101111",
      "010110000000000000000111100011111110101011011101111000011010100111110010101100101110010" when "010110000",
      "010110001000000000000111101001011111101011000001101011110010001000111101001011110011000" when "010110001",
      "010110010000000000000111101111000010101010100101100001111010101001111010100010011011111" when "010110010",
      "010110011000000000000111110100100111101010001001011010110101001010101010110010101101110" when "010110011",
      "010110100000000000000111111010001110101001101101010110100010101011001101111110101110101" when "010110100",
      "010110101000000000000111111111110111101001010001010101000100001011100100001000100101001" when "010110101",
      "010110110000000000001000000101100010101000110101010110011010101011101101010010011000100" when "010110110",
      "010110111000000000001000001011001111101000011001011010100111001011101001011110010001000" when "010110111",
      "010111000000000000001000010000111110100111111101100001101010101011011000101110010111100" when "010111000",
      "010111001000000000001000010110101111100111100001101011100110001010111011000100110101011" when "010111001",
      "010111010000000000001000011100100010100111000101111000011010101010010000100011110101010" when "010111010",
      "010111011000000000001000100010010111100110101010001000001001001001011001001101100010010" when "010111011",
      "010111100000000000001000101000001110100110001110011010110010101000010101000100001000010" when "010111100",
      "010111101000000000001000101110000111100101110010110000011000000111000100001001110011110" when "010111101",
      "010111110000000000001000110100000010100101010111001000111010100101100110100000110010010" when "010111110",
      "010111111000000000001000111001111111100100111011100100011011000011111100001011010001110" when "010111111",
      "011000000000000000001000111111111110100100100000000010111010100010000101001011100001001" when "011000000",
      "011000001000000000001001000101111111100100000100100100011010000000000001100011110000001" when "011000001",
      "011000010000000000001001001100000010100011101001001000111010011101110001010110001111000" when "011000010",
      "011000011000000000001001010010000111100011001101110000011100111011010100100101001111000" when "011000011",
      "011000100000000000001001011000001110100010110010011011000010011000101011010011000001110" when "011000100",
      "011000101000000000001001011110010111100010010111001000101011110101110101100001111010010" when "011000101",
      "011000110000000000001001100100100010100001111011111001011010010010110011010100001011100" when "011000110",
      "011000111000000000001001101010101111100001100000101101001110101111100100101100001010000" when "011000111",
      "011001000000000000001001110000111110100001000101100100001010001100001001101100001010010" when "011001000",
      "011001001000000000001001110111001111100000101010011110001101101000100010010110100010000" when "011001001",
      "011001010000000000001001111101100010100000001111011011011010000100101110101101100111110" when "011001010",
      "011001011000000000001010000011110111011111110100011011110000100000101110110011110010100" when "011001011",
      "011001100000000000001010001010001110011111011001011111010001111100100010101011011010010" when "011001100",
      "011001101000000000001010010000100111011110111110100101111111011000001010010110110111100" when "011001101",
      "011001110000000000001010010111000010011110100011101111111001110011100101111000100011100" when "011001110",
      "011001111000000000001010011101011111011110001000111101000010001110110101010010111000101" when "011001111",
      "011010000000000000001010100011111110011101101110001101011001101001111000101000010001101" when "011010000",
      "011010001000000000001010101010011111011101010011100001000001000100101111111011001010010" when "011010001",
      "011010010000000000001010110001000010011100111000110111111001011111011011001101111110101" when "011010010",
      "011010011000000000001010110111100111011100011110010010000011111001111010100011001100000" when "011010011",
      "011010100000000000001010111110001110011100000011101111100001010100001101111101010000011" when "011010100",
      "011010101000000000001011000100110111011011101001010000010010101110010101011110101010010" when "011010101",
      "011010110000000000001011001011100010011011001110110100011001001000010001001001111001000" when "011010110",
      "011010111000000000001011010010001111011010110100011011110101100010000001000001011100110" when "011010111",
      "011011000000000000001011011000111110011010011010000110101000111011100101000111110110011" when "011011000",
      "011011001000000000001011011111101111011001111111110100110100010100111101011111100111100" when "011011001",
      "011011010000000000001011100110100010011001100101100110011000101110001010001011010010100" when "011011010",
      "011011011000000000001011101101010111011001001011011011010111000111001011001101011010100" when "011011011",
      "011011100000000000001011110100001110011000110001010011110000100000000000101000100011011" when "011011100",
      "011011101000000000001011111011000111011000010111001111100101111000101010011111010001110" when "011011101",
      "011011110000000000001100000010000010010111111101001110111000010001001000110100001011000" when "011011110",
      "011011111000000000001100001000111111010111100011010001101000101001011011101001110101010" when "011011111",
      "011100000000000000001100001111111110010111001001010111111000000001100011000010110111011" when "011100000",
      "011100001000000000001100010110111111010110101111100001100111011001011111000001111001000" when "011100001",
      "011100010000000000001100011110000010010110010101101110110111110001001111101001100010100" when "011100010",
      "011100011000000000001100100101000111010101111011111111101010001000110100111100011100111" when "011100011",
      "011100100000000000001100101100001110010101100010010011111111100000001110111101010010010" when "011100100",
      "011100101000000000001100110011010111010101001000101011111000110111011101101110101101000" when "011100101",
      "011100110000000000001100111010100010010100101111000111010111001110100001010011011000101" when "011100110",
      "011100111000000000001101000001101111010100010101100110011011100101011001101110000001010" when "011100111",
      "011101000000000000001101001000111110010011111100001001000110111100000111000001010011110" when "011101000",
      "011101001000000000001101010000001111010011100010101111011010010010101001001111111101110" when "011101001",
      "011101010000000000001101010111100010010011001001011001010110101001000000011100101101100" when "011101010",
      "011101011000000000001101011110110111010010110000000110111100111111001100101010010010010" when "011101011",
      "011101100000000000001101100110001110010010010110111000001110010101001101111011011100000" when "011101100",
      "011101101000000000001101101101100111010001111101101101001011101011000100010010111011000" when "011101101",
      "011101110000000000001101110101000010010001100100100101110110000000101111110011100001000" when "011101110",
      "011101111000000000001101111100011111010001001011100010001110010110010000011111111111111" when "011101111",
      "011110000000000000001110000011111110010000110010100010010101101011100110011011001010101" when "011110000",
      "011110001000000000001110001011011111010000011001100110001101000000110001100111110100110" when "011110001",
      "011110010000000000001110010011000010010000000000101101110101010101110010001000110010111" when "011110010",
      "011110011000000000001110011010100111001111100111111001001111101010101000000000111001111" when "011110011",
      "011110100000000000001110100010001110001111001111001000011100111111010011010010111111110" when "011110100",
      "011110101000000000001110101001110111001110110110011011011110010011110100000001111011000" when "011110101",
      "011110110000000000001110110001100010001110011101110010010100101000001010010000100011000" when "011110110",
      "011110111000000000001110111001001111001110000101001101000000111100010110000001110000001" when "011110111",
      "011111000000000000001111000000111110001101101100101011100100010000010111011000011011000" when "011111000",
      "011111001000000000001111001000101111001101010100001101111111100100001110010111011101011" when "011111001",
      "011111010000000000001111010000100010001100111011110100010011110111111011000001110001100" when "011111010",
      "011111011000000000001111011000010111001100100011011110100010001011011101011010010010110" when "011111011",
      "011111100000000000001111100000001110001100001011001100101011011110110101100011111100101" when "011111100",
      "011111101000000000001111101000000111001011110010111110110000110010000011100001101100000" when "011111101",
      "011111110000000000001111110000000010001011011010110100110011000101000111010110011110010" when "011111110",
      "011111111000000000001111110111111111001011000010101110110011011000000001000101010001010" when "011111111",
      "100000000000000000001111111111111110001010101010101100110010101010110000110001000100010" when "100000000",
      "100000001000000000010000000111111111001010010010101110110001111101010110011100110110101" when "100000001",
      "100000010000000000010000010000000010001001111010110100110010001111110010001011101000111" when "100000010",
      "100000011000000000010000011000000111001001100010111110110100100010000100000000011100000" when "100000011",
      "100000100000000000010000100000001110001001001011001100111001110100001011111110010001111" when "100000100",
      "100000101000000000010000101000010111001000110011011111000011000110001010001000001101010" when "100000101",
      "100000110000000000010000110000100010001000011011110101010001010111111110100001010001100" when "100000110",
      "100000111000000000010000111000101111001000000100001111100101101001101001001100100010101" when "100000111",
      "100001000000000000010001000000111110000111101100101110000000111011001010001101000101100" when "100001000",
      "100001001000000000010001001001001111000111010101010000100100001100100001100101111111110" when "100001001",
      "100001010000000000010001010001100010000110111101110111010000011101101111011010011000000" when "100001010",
      "100001011000000000010001011001110111000110100110100010000110101110110011101101010101000" when "100001011",
      "100001100000000000010001100010001110000110001111010001000111111111101110100001111110111" when "100001100",
      "100001101000000000010001101010100111000101111000000100010101010000011111111011011110001" when "100001101",
      "100001110000000000010001110011000010000101100000111011101111100001000111111100111100010" when "100001110",
      "100001111000000000010001111011011111000101001001110111010111110001100110101001100011010" when "100001111",
      "100010000000000000010010000011111110000100110010110111001111000001111100000100011110000" when "100010000",
      "100010001000000000010010001100011111000100011011111011010110010010001000010000111000001" when "100010001",
      "100010010000000000010010010101000010000100000101000011101110100010001011010001111110001" when "100010010",
      "100010011000000000010010011101100111000011101110010000011000110010000101001010111101000" when "100010011",
      "100010100000000000010010100110001110000011010111100001010110000001110101111111000010110" when "100010100",
      "100010101000000000010010101110110111000011000000110110100111010001011101110001011101111" when "100010101",
      "100010110000000000010010110111100010000010101010010000001101100000111100100101011101110" when "100010110",
      "100010111000000000010011000000001111000010010011101110001001110000010010011110010010100" when "100010111",
      "100011000000000000010011001000111110000001111101010000011100111111011111011111001101001" when "100011000",
      "100011001000000000010011010001101111000001100110110111001000001110100011101011011111000" when "100011001",
      "100011010000000000010011011010100010000001010000100010001100011101011111000110011010110" when "100011010",
      "100011011000000000010011100011010111000000111010010001101010101100010001110011010011100" when "100011011",
      "100011100000000000010011101100001110000000100100000101100011111010111011110101011100111" when "100011100",
      "100011101000000000010011110101000111000000001101111101111001001001011101010000001011110" when "100011101",
      "100011110000000000010011111110000001111111110111111010101011010111110110000110110101011" when "100011110",
      "100011111000000000010100000110111110111111100001111011111011100110000110011100101111111" when "100011111",
      "100100000000000000010100001111111101111111001100000001101010110100001110010101010010001" when "100100000",
      "100100001000000000010100011000111110111110110110001011111010000010001101110011110011111" when "100100001",
      "100100010000000000010100100010000001111110100000011010101010010000000100111011101101010" when "100100010",
      "100100011000000000010100101011000110111110001010101101111100011101110011110000010111101" when "100100011",
      "100100100000000000010100110100001101111101110101000101110001101011011010010101001100110" when "100100100",
      "100100101000000000010100111101010110111101011111100010001010111000111000101101100111010" when "100100101",
      "100100110000000000010101000110100001111101001010000011001001000110001110111101000010100" when "100100110",
      "100100111000000000010101001111101110111100110100101000101101010011011101000110111010101" when "100100111",
      "100101000000000000010101011000111101111100011111010010111000100000100011001110101100101" when "100101000",
      "100101001000000000010101100010001110111100001010000001101011101101100001010111110101111" when "100101001",
      "100101010000000000010101101011100001111011110100110101000111111010010111100101110101000" when "100101010",
      "100101011000000000010101110100110110111011011111101101001110000111000101111100001001000" when "100101011",
      "100101100000000000010101111110001101111011001010101001111111010011101100011110010001101" when "100101100",
      "100101101000000000010110000111100110111010110101101011011100100000001011001111101111110" when "100101101",
      "100101110000000000010110010001000001111010100000110001100110101100100010010100000100101" when "100101110",
      "100101111000000000010110011010011110111010001011111100011110111000110001101110110010011" when "100101111",
      "100110000000000000010110100011111101111001110111001100000110000100111001100011011011111" when "100110000",
      "100110001000000000010110101101011110111001100010100000011101010000111001110101100100111" when "100110001",
      "100110010000000000010110110111000001111001001101111001100101011100110010101000110001100" when "100110010",
      "100110011000000000010111000000100110111000111001010111011111101000100100000000100111000" when "100110011",
      "100110100000000000010111001010001101111000100100111010001100110100001110000000101011010" when "100110100",
      "100110101000000000010111010011110110111000010000100001101101111111110000101100100100111" when "100110101",
      "100110110000000000010111011101100001110111111100001110000100001011001100000111111011011" when "100110110",
      "100110111000000000010111100111001110110111100111111111010000010110100000010110010110101" when "100110111",
      "100111000000000000010111110000111101110111010011110101010011100001101101011011011111101" when "100111000",
      "100111001000000000010111111010101110110110111111110000001110101100110011011011000000001" when "100111001",
      "100111010000000000011000000100100001110110101011110000000010110111110010011000100010010" when "100111010",
      "100111011000000000011000001110010110110110010111110100110001000010101010010111110001010" when "100111011",
      "100111100000000000011000011000001101110110000011111110011010001101011011011100011001000" when "100111100",
      "100111101000000000011000100010000110110101110000001100111111011000000101101010000110010" when "100111101",
      "100111110000000000011000101100000001110101011100100000100001100010101001000100100110001" when "100111110",
      "100111111000000000011000110101111110110101001000111001000001101101000101101111100110111" when "100111111",
      "101000000000000000011000111111111101110100110101010110100000110111011011101110110111011" when "101000000",
      "101000001000000000011001001001111110110100100001111001000000000001101011000110000111010" when "101000001",
      "101000010000000000011001010100000001110100001110100000100000001011110011111001000110111" when "101000010",
      "101000011000000000011001011110000110110011111011001101000010010101110110001011100111011" when "101000011",
      "101000100000000000011001101000001101110011100111111110100111011111110010000001011010101" when "101000100",
      "101000101000000000011001110010010110110011010100110101010000101001100111011110010011010" when "101000101",
      "101000110000000000011001111100100001110011000001110000111110110011010110100110000100101" when "101000110",
      "101000111000000000011010000110101110110010101110110001110010111100111111011100100010110" when "101000111",
      "101001000000000000011010010000111101110010011011110111101110000110100010000101100010110" when "101001000",
      "101001001000000000011010011011001110110010001001000010110001001111111110100100111010000" when "101001001",
      "101001010000000000011010100101100001110001110110010010111101011001010100111110011111001" when "101001010",
      "101001011000000000011010101111110110110001100011101000010011100010100101010110001001000" when "101001011",
      "101001100000000000011010111010001101110001010001000010110100101011101111101111101111101" when "101001100",
      "101001101000000000011011000100100110110000111110100010100001110100110100001111001011110" when "101001101",
      "101001110000000000011011001111000001110000101100000111011011111101110010111000010110100" when "101001110",
      "101001111000000000011011011001011110110000011001110001100100000110101011101111001010001" when "101001111",
      "101010000000000000011011100011111101110000000111100000111011001111011110110111100001011" when "101010000",
      "101010001000000000011011101110011110101111110101010101100010011000001100010101011000001" when "101010001",
      "101010010000000000011011111001000001101111100011001111011010100000110100001100101010101" when "101010010",
      "101010011000000000011100000011100110101111010001001110100100101001010110100001010101111" when "101010011",
      "101010100000000000011100001110001101101110111111010011000001110001110011010111010111111" when "101010100",
      "101010101000000000011100011000110110101110101101011100110010111010001010110010101111011" when "101010101",
      "101010110000000000011100100011100001101110011011101011111001000010011100110111011011100" when "101010110",
      "101010111000000000011100101110001110101110001010000000010101001010101001101001011100100" when "101010111",
      "101011000000000000011100111000111101101101111000011010001000010010110001001100110011010" when "101011000",
      "101011001000000000011101000011101110101101100110111001010011011010110011100101100001010" when "101011001",
      "101011010000000000011101001110100001101101010101011101110111100010110000110111101001001" when "101011010",
      "101011011000000000011101011001010110101101000100000111110101101010101001000111001101110" when "101011011",
      "101011100000000000011101100100001101101100110010110111001110110010011100011000010011001" when "101011100",
      "101011101000000000011101101111000110101100100001101100000011111010001010101110111110000" when "101011101",
      "101011110000000000011101111010000001101100010000100110010110000001110100001111010011100" when "101011110",
      "101011111000000000011110000100111110101011111111100110000110001001011000111101011001110" when "101011111",
      "101100000000000000011110001111111101101011101110101011010101010000111000111101010111111" when "101100000",
      "101100001000000000011110011010111110101011011101110110000100011000010100010011010101011" when "101100001",
      "101100010000000000011110100110000001101011001101000110010100011111101011000011011010100" when "101100010",
      "101100011000000000011110110001000110101010111100011100000110100110111101010001110000100" when "101100011",
      "101100100000000000011110111100001101101010101011110111011011101110001011000010100001010" when "101100100",
      "101100101000000000011111000111010110101010011011011000010100110101010100011001110111011" when "101100101",
      "101100110000000000011111010010100001101010001010111110110010111100011001011011111110010" when "101100110",
      "101100111000000000011111011101101110101001111010101010110111000011011010001101000010000" when "101100111",
      "101101000000000000011111101000111101101001101010011100100010001010010110110001001111011" when "101101000",
      "101101001000000000011111110100001110101001011010010011110101010001001111001100110100001" when "101101001",
      "101101010000000000011111111111100001101001001010010000110001011000000011100011111110101" when "101101010",
      "101101011000000000100000001010110110101000111010010011010111011110110011111010111110000" when "101101011",
      "101101100000000000100000010110001101101000101010011011101000100101100000010110000010001" when "101101100",
      "101101101000000000100000100001100110101000011010101001100101101100001000111001011011101" when "101101101",
      "101101110000000000100000101101000001101000001010111101001111110010101101101001011011110" when "101101110",
      "101101111000000000100000111000011110100111111011010110100111111001001110101010010100111" when "101101111",
      "101110000000000000100001000011111101100111101011110101101110111111101100000000011001101" when "101110000",
      "101110001000000000100001001111011110100111011100011010100110000110000101101111111101110" when "101110001",
      "101110010000000000100001011011000001100111001101000101001110001100011011111101010101101" when "101110010",
      "101110011000000000100001100110100110100110111101110101101000010010101110101100110110011" when "101110011",
      "101110100000000000100001110010001101100110101110101011110101011000111110000010110101110" when "101110100",
      "101110101000000000100001111101110110100110011111100111110110011111001010000011101010101" when "101110101",
      "101110110000000000100010001001100001100110010000101001101100100101010010110011101100001" when "101110110",
      "101110111000000000100010010101001110100110000001110001011000101011011000010111010010100" when "101110111",
      "101111000000000000100010100000111101100101110010111110111011110001011010110010110110101" when "101111000",
      "101111001000000000100010101100101110100101100100010010010110110111011010001010110010001" when "101111001",
      "101111010000000000100010111000100001100101010101101011101010111101010110100011011111011" when "101111010",
      "101111011000000000100011000100010110100101000111001010111001000011010000000001011001011" when "101111011",
      "101111100000000000100011010000001101100100111000110000000010001001000110101000111100010" when "101111100",
      "101111101000000000100011011100000110100100101010011011000111001110111010011110100100011" when "101111101",
      "101111110000000000100011101000000001100100011100001100001001010100101011100110101111010" when "101111110",
      "101111111000000000100011110011111110100100001110000011001001011010011010000101111011000" when "101111111",
      "110000000000000000100011111111111101100100000000000000001000100000000110000000100110100" when "110000000",
      "110000001000000000100100001011111110100011110010000011000111100101101111011011010001011" when "110000001",
      "110000010000000000100100011000000001100011100100001100000111101011010110011010011100000" when "110000010",
      "110000011000000000100100100100000110100011010110011011001001110000111011000010100111011" when "110000011",
      "110000100000000000100100110000001101100011001000110000001110110110011101011000010101100" when "110000100",
      "110000101000000000100100111100010110100010111011001011010111111011111101100000001001001" when "110000101",
      "110000110000000000100101001000100001100010101101101100100110000001011011011110100101011" when "110000110",
      "110000111000000000100101010100101110100010100000010011111010000110110111011000001110100" when "110000111",
      "110001000000000000100101100000111101100010010011000001010101001100010001010001101001011" when "110001000",
      "110001001000000000100101101101001110100010000101110100111000010001101001001111011011101" when "110001001",
      "110001010000000000100101111001100001100001111000101110100100010110111111010110001011101" when "110001010",
      "110001011000000000100110000101110110100001101011101110011010011100010011101010100000011" when "110001011",
      "110001100000000000100110010010001101100001011110110100011011100001100110010001000010000" when "110001100",
      "110001101000000000100110011110100110100001010010000000101000100110110111001110011001000" when "110001101",
      "110001110000000000100110101011000001100001000101010011000010101100000110100111001110101" when "110001110",
      "110001111000000000100110110111011110100000111000101011101010110001010100100000001101010" when "110001111",
      "110010000000000000100111000011111101100000101100001010100001110110100000111101111111100" when "110010000",
      "110010001000000000100111010000011110100000011111101111101000111011101100000101010001001" when "110010001",
      "110010010000000000100111011101000001100000010011011011000001000000110101111010101110100" when "110010010",
      "110010011000000000100111101001100110100000000111001100101011000101111110100011000100111" when "110010011",
      "110010100000000000100111110110001101011111111011000100101000001011000110000011000001111" when "110010100",
      "110010101000000000101000000010110110011111101111000010111001010000001100011111010100010" when "110010101",
      "110010110000000000101000001111100001011111100011000111011111010101010001111100101011011" when "110010110",
      "110010111000000000101000011100001110011111010111010010011011011010010110011111110111011" when "110010111",
      "110011000000000000101000101000111101011111001011100011101110011111011010001101101001001" when "110011000",
      "110011001000000000101000110101101110011110111111111011011001100100011101001010110010010" when "110011001",
      "110011010000000000101001000010100001011110110100011001011101101001011111011100000101001" when "110011010",
      "110011011000000000101001001111010110011110101000111101111011101110100001000110010100111" when "110011011",
      "110011100000000000101001011100001101011110011101101000110100110011100010001110010101011" when "110011100",
      "110011101000000000101001101001000110011110010010011010001001111000100010111000111011010" when "110011101",
      "110011110000000000101001110110000001011110000111010001111011111101100011001010111011111" when "110011110",
      "110011111000000000101010000010111110011101111100010000001100000010100011001001001101011" when "110011111",
      "110100000000000000101010001111111101011101110001010100111011000111100010111000100110101" when "110100000",
      "110100001000000000101010011100111110011101100110100000001010001100100010011101111111010" when "110100001",
      "110100010000000000101010101010000001011101011011110001111010010001100001111110001111101" when "110100010",
      "110100011000000000101010110111000110011101010001001010001100010110100001011110010001000" when "110100011",
      "110100100000000000101011000100001101011101000110101001000001011011100001000010111101000" when "110100100",
      "110100101000000000101011010001010110011100111100001110011010100000100000110001001110011" when "110100101",
      "110100110000000000101011011110100001011100110001111010011000100101100000101110000000101" when "110100110",
      "110100111000000000101011101011101110011100100111101100111100101010100000111110001111101" when "110100111",
      "110101000000000000101011111000111101011100011101100110000111101111100001100110111000100" when "110101000",
      "110101001000000000101100000110001110011100010011100101111010110100100010101100111000110" when "110101001",
      "110101010000000000101100010011100001011100001001101100010110111001100100010101001110101" when "110101010",
      "110101011000000000101100100000110110011011111111111001011100111110100110100100111001100" when "110101011",
      "110101100000000000101100101110001101011011110110001101001110000011101001100000111001010" when "110101100",
      "110101101000000000101100111011100110011011101100100111101011001000101101001110001110010" when "110101101",
      "110101110000000000101101001001000001011011100011001000110101001101110001110001111010000" when "110101110",
      "110101111000000000101101010110011110011011011001110000101101010010110111010000111110110" when "110101111",
      "110110000000000000101101100011111101011011010000011111010100010111111101110000011111001" when "110110000",
      "110110001000000000101101110001011110011011000111010100101011011101000101010101011111000" when "110110001",
      "110110010000000000101101111111000001011010111110010000110011100010001110000101000010110" when "110110010",
      "110110011000000000101110001100100110011010110101010011101101100111011000000100001111010" when "110110011",
      "110110100000000000101110011010001101011010101100011101011010101100100011011000001010100" when "110110100",
      "110110101000000000101110100111110110011010100011101101111011110001110000000101111011010" when "110110101",
      "110110110000000000101110110101100001011010011011000101010001110110111110010010101000110" when "110110110",
      "110110111000000000101111000011001110011010010010100011011101111100001110000011011011001" when "110110111",
      "110111000000000000101111010000111101011010001010001000100001000001011111011101011011011" when "110111000",
      "110111001000000000101111011110101110011010000001110100011100000110110010100101110010111" when "110111001",
      "110111010000000000101111101100100001011001111001100111010000001100000111100001101100010" when "110111010",
      "110111011000000000101111111010010110011001110001100000111110010001011110010110010010101" when "110111011",
      "110111100000000000110000001000001101011001101001100001100111010110110111001000110001101" when "110111100",
      "110111101000000000110000010110000110011001100001101001001100011100010001111110010110001" when "110111101",
      "110111110000000000110000100100000001011001011001110111101110100001101110111100001101011" when "110111110",
      "110111111000000000110000110001111110011001010010001101001110100111001110000111100101101" when "110111111",
      "111000000000000000110000111111111101011001001010101001101101101100101111100101101101101" when "111000000",
      "111000001000000000110001001101111110011001000011001101001100110010010011011011110101000" when "111000001",
      "111000010000000000110001011100000001011000111011110111101100110111111001101111001100010" when "111000010",
      "111000011000000000110001101010000110011000110100101001001110111101100010100101000100011" when "111000011",
      "111000100000000000110001111000001101011000101101100001110100000011001110000010101111010" when "111000100",
      "111000101000000000110010000110010110011000100110100001011101001000111100001101011111101" when "111000101",
      "111000110000000000110010010100100001011000011111101000001011001110101101001010101000110" when "111000110",
      "111000111000000000110010100010101110011000011000110101111111010100100000111111011110111" when "111000111",
      "111001000000000000110010110000111101011000010010001010111010011010010111110001010110110" when "111001000",
      "111001001000000000110010111111001110011000001011100110111101100000010001100101100110001" when "111001001",
      "111001010000000000110011001101100001011000000101001010001001100110001110100001100011010" when "111001010",
      "111001011000000000110011011011110110010111111110110100011111101100001110101010100101011" when "111001011",
      "111001100000000000110011101010001101010111111000100110000000110010010010000110000100010" when "111001100",
      "111001101000000000110011111000100110010111110010011110101101111000011000111001011000100" when "111001101",
      "111001110000000000110100000111000001010111101100011110100111111110100011001001111011101" when "111001110",
      "111001111000000000110100010101011110010111100110100101110000000100110000111101000111110" when "111001111",
      "111010000000000000110100100011111101010111100000110100000111001011000010011000010111101" when "111010000",
      "111010001000000000110100110010011110010111011011001001101110010001010111100001000111000" when "111010001",
      "111010010000000000110101000001000001010111010101100110100110010111110000011100110010010" when "111010010",
      "111010011000000000110101001111100110010111010000001010110000011110001101010000110110011" when "111010011",
      "111010100000000000110101011110001101010111001010110110001101100100101110000010110001010" when "111010100",
      "111010101000000000110101101100110110010111000101101000111110101011010010111000000001110" when "111010101",
      "111010110000000000110101111011100001010111000000100011000100110001111011110110000110111" when "111010110",
      "111010111000000000110110001010001110010110111011100100100000111000101001000010100001001" when "111010111",
      "111011000000000000110110011000111101010110110110101101010011111111011010100010110001001" when "111011000",
      "111011001000000000110110100111101110010110110001111101011111000110010000011100011000101" when "111011001",
      "111011010000000000110110110110100001010110101101010101000011001101001010110100111010000" when "111011010",
      "111011011000000000110111000101010110010110101000110100000001010100001001110001111000011" when "111011011",
      "111011100000000000110111010100001101010110100100011010011010011011001101011000110111100" when "111011100",
      "111011101000000000110111100011000110010110100000001000001111100010010101101111011100001" when "111011101",
      "111011110000000000110111110010000001010110011011111101100001101001100010111011001011101" when "111011110",
      "111011111000000000111000000000111110010110010111111010010001110000110101000001101100000" when "111011111",
      "111100000000000000111000001111111101010110010011111110100000111000001100001000100100011" when "111100000",
      "111100001000000000111000011110111110010110010000001010001111111111101000010101011100001" when "111100001",
      "111100010000000000111000101110000001010110001100011101100000000111001001101101111011110" when "111100010",
      "111100011000000000111000111101000110010110001000111000010010001110110000010111101100011" when "111100011",
      "111100100000000000111001001100001101010110000101011010100111010110011100011000010111111" when "111100100",
      "111100101000000000111001011011010110010110000010000100100000011110001101110101101000111" when "111100101",
      "111100110000000000111001101010100001010101111110110101111110100110000100110101001010110" when "111100110",
      "111100111000000000111001111001101110010101111011101111000010101110000001011100101001100" when "111100111",
      "111101000000000000111010001000111101010101111000101111101101110110000011110001110010010" when "111101000",
      "111101001000000000111010011000001110010101110101111000000000111110001011111010010010100" when "111101001",
      "111101010000000000111010100111100001010101110011000111111101000110011001111011111000100" when "111101010",
      "111101011000000000111010110110110110010101110000011111100011001110101101111100010011101" when "111101011",
      "111101100000000000111011000110001101010101101101111110110100010111001000000001010011101" when "111101100",
      "111101101000000000111011010101100110010101101011100101110001011111101000010000101001001" when "111101101",
      "111101110000000000111011100101000001010101101001010100011011101000001110110000000101100" when "111101110",
      "111101111000000000111011110100011110010101100111001010110011110000111011100101011010111" when "111101111",
      "111110000000000000111100000011111101010101100101001000111010111001101110110110011100001" when "111110000",
      "111110001000000000111100010011011110010101100011001110110010000010101000101000111100111" when "111110001",
      "111110010000000000111100100011000001010101100001011100011010001011101001000010110001101" when "111110010",
      "111110011000000000111100110010100110010101011111110001110100010100110000001001101111010" when "111110011",
      "111110100000000000111101000010001101010101011110001111000001011101111110000011101011111" when "111110100",
      "111110101000000000111101010001110110010101011100110100000010100111010010110110011110000" when "111110101",
      "111110110000000000111101100001100001010101011011100000111000110000101110100111111101000" when "111110110",
      "111110111000000000111101110001001110010101011010010101100100111010010001011110000001001" when "111110111",
      "111111000000000000111110000000111101010101011001010010001000000011111011011110100011001" when "111111000",
      "111111001000000000111110010000101110010101011000010110100011001101101100101111011100101" when "111111001",
      "111111010000000000111110100000100001010101010111100010110111010111100101010110101000001" when "111111010",
      "111111011000000000111110110000010110010101010110110111000101100001100101011010000000101" when "111111011",
      "111111100000000000111111000000001101010101010110010011001110101011101100111111100010000" when "111111100",
      "111111101000000000111111010000000110010101010101110111010011110101111100001101001001000" when "111111101",
      "111111110000000000111111100000000001010101010101100011010110000000010011001000110010111" when "111111110",
      "111111111000000000111111101111111110010101010101010111010110001010110001111000011101111" when "111111111",
      "---------------------------------------------------------------------------------------" when others;
   Y1_c4 <= Y0_c4; -- for the possible blockram register
   Y <= Y1_c4;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_104_Freq300_uid48
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_104_Freq300_uid48 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(103 downto 0);
          Y : in  std_logic_vector(103 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(103 downto 0)   );
end entity;

architecture arch of IntAdder_104_Freq300_uid48 is
signal Rtmp_c4 :  std_logic_vector(103 downto 0);
signal X_c3, X_c4 :  std_logic_vector(103 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               X_c3 <= X;
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               X_c4 <= X_c3;
               Cin_c4 <= Cin_c3;
            end if;
         end if;
      end process;
   Rtmp_c4 <= X_c4 + Y + Cin_c4;
   R <= Rtmp_c4;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable3_Freq300_uid50
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable3_Freq300_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(78 downto 0)   );
end entity;

architecture arch of LogTable3_Freq300_uid50 is
signal Y0_c5 :  std_logic_vector(78 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c5 :  std_logic_vector(78 downto 0);
begin
   with X  select  Y0_c5 <= 
      "0000000000000000000000000000000000000000000000000000000000000000000000000001000" when "0000000000",
      "0000000001000000000000000000000000000000000000111111111111110000000000000001000" when "0000000001",
      "0000000010000000000000000000000000000000000011111111111111100000000000000001001" when "0000000010",
      "0000000011000000000000000000000000000000001000111111111111010000000000000001100" when "0000000011",
      "0000000100000000000000000000000000000000001111111111111111000000000000000010011" when "0000000100",
      "0000000101000000000000000000000000000000011000111111111110110000000000000011101" when "0000000101",
      "0000000110000000000000000000000000000000100011111111111110100000000000000101100" when "0000000110",
      "0000000111000000000000000000000000000000110000111111111110010000000000001000001" when "0000000111",
      "0000001000000000000000000000000000000000111111111111111110000000000000001011101" when "0000001000",
      "0000001001000000000000000000000000000001010000111111111101110000000000010000010" when "0000001001",
      "0000001010000000000000000000000000000001100011111111111101100000000000010101111" when "0000001010",
      "0000001011000000000000000000000000000001111000111111111101010000000000011100110" when "0000001011",
      "0000001100000000000000000000000000000010001111111111111101000000000000100101000" when "0000001100",
      "0000001101000000000000000000000000000010101000111111111100110000000000101110110" when "0000001101",
      "0000001110000000000000000000000000000011000011111111111100100000000000111010001" when "0000001110",
      "0000001111000000000000000000000000000011100000111111111100010000000001000111010" when "0000001111",
      "0000010000000000000000000000000000000011111111111111111100000000000001010110011" when "0000010000",
      "0000010001000000000000000000000000000100100000111111111011110000000001100111011" when "0000010001",
      "0000010010000000000000000000000000000101000011111111111011100000000001111010100" when "0000010010",
      "0000010011000000000000000000000000000101101000111111111011010000000010001111111" when "0000010011",
      "0000010100000000000000000000000000000110001111111111111011000000000010100111101" when "0000010100",
      "0000010101000000000000000000000000000110111000111111111010110000000011000010000" when "0000010101",
      "0000010110000000000000000000000000000111100011111111111010100000000011011110111" when "0000010110",
      "0000010111000000000000000000000000001000010000111111111010010000000011111110100" when "0000010111",
      "0000011000000000000000000000000000001000111111111111111010000000000100100001000" when "0000011000",
      "0000011001000000000000000000000000001001110000111111111001110000000101000110100" when "0000011001",
      "0000011010000000000000000000000000001010100011111111111001100000000101101111001" when "0000011010",
      "0000011011000000000000000000000000001011011000111111111001010000000110011011000" when "0000011011",
      "0000011100000000000000000000000000001100001111111111111001000000000111001010011" when "0000011100",
      "0000011101000000000000000000000000001101001000111111111000110000000111111101001" when "0000011101",
      "0000011110000000000000000000000000001110000011111111111000100000001000110011100" when "0000011110",
      "0000011111000000000000000000000000001111000000111111111000010000001001101101101" when "0000011111",
      "0000100000000000000000000000000000001111111111111111111000000000001010101011101" when "0000100000",
      "0000100001000000000000000000000000010001000000111111110111110000001011101101110" when "0000100001",
      "0000100010000000000000000000000000010010000011111111110111100000001100110011111" when "0000100010",
      "0000100011000000000000000000000000010011001000111111110111010000001101111110010" when "0000100011",
      "0000100100000000000000000000000000010100001111111111110111000000001111001101000" when "0000100100",
      "0000100101000000000000000000000000010101011000111111110110110000010000100000010" when "0000100101",
      "0000100110000000000000000000000000010110100011111111110110100000010001111000001" when "0000100110",
      "0000100111000000000000000000000000010111110000111111110110010000010011010100110" when "0000100111",
      "0000101000000000000000000000000000011000111111111111110110000000010100110110011" when "0000101000",
      "0000101001000000000000000000000000011010010000111111110101110000010110011100111" when "0000101001",
      "0000101010000000000000000000000000011011100011111111110101100000011000001000100" when "0000101010",
      "0000101011000000000000000000000000011100111000111111110101010000011001111001011" when "0000101011",
      "0000101100000000000000000000000000011110001111111111110101000000011011101111101" when "0000101100",
      "0000101101000000000000000000000000011111101000111111110100110000011101101011100" when "0000101101",
      "0000101110000000000000000000000000100001000011111111110100100000011111101100111" when "0000101110",
      "0000101111000000000000000000000000100010100000111111110100010000100001110100000" when "0000101111",
      "0000110000000000000000000000000000100011111111111111110100000000100100000001000" when "0000110000",
      "0000110001000000000000000000000000100101100000111111110011110000100110010100000" when "0000110001",
      "0000110010000000000000000000000000100111000011111111110011100000101000101101001" when "0000110010",
      "0000110011000000000000000000000000101000101000111111110011010000101011001100100" when "0000110011",
      "0000110100000000000000000000000000101010001111111111110011000000101101110010011" when "0000110100",
      "0000110101000000000000000000000000101011111000111111110010110000110000011110101" when "0000110101",
      "0000110110000000000000000000000000101101100011111111110010100000110011010001100" when "0000110110",
      "0000110111000000000000000000000000101111010000111111110010010000110110001011001" when "0000110111",
      "0000111000000000000000000000000000110000111111111111110010000000111001001011101" when "0000111000",
      "0000111001000000000000000000000000110010110000111111110001110000111100010011001" when "0000111001",
      "0000111010000000000000000000000000110100100011111111110001100000111111100001111" when "0000111010",
      "0000111011000000000000000000000000110110011000111111110001010001000010110111110" when "0000111011",
      "0000111100000000000000000000000000111000001111111111110001000001000110010101000" when "0000111100",
      "0000111101000000000000000000000000111010001000111111110000110001001001111001110" when "0000111101",
      "0000111110000000000000000000000000111100000011111111110000100001001101100110001" when "0000111110",
      "0000111111000000000000000000000000111110000000111111110000010001010001011010010" when "0000111111",
      "0001000000000000000000000000000000111111111111111111110000000001010101010110011" when "0001000000",
      "0001000001000000000000000000000001000010000000111111101111110001011001011010011" when "0001000001",
      "0001000010000000000000000000000001000100000011111111101111100001011101100110100" when "0001000010",
      "0001000011000000000000000000000001000110001000111111101111010001100001111010111" when "0001000011",
      "0001000100000000000000000000000001001000001111111111101111000001100110010111101" when "0001000100",
      "0001000101000000000000000000000001001010011000111111101110110001101010111100111" when "0001000101",
      "0001000110000000000000000000000001001100100011111111101110100001101111101010111" when "0001000110",
      "0001000111000000000000000000000001001110110000111111101110010001110100100001100" when "0001000111",
      "0001001000000000000000000000000001010000111111111111101110000001111001100001000" when "0001001000",
      "0001001001000000000000000000000001010011010000111111101101110001111110101001100" when "0001001001",
      "0001001010000000000000000000000001010101100011111111101101100010000011111011001" when "0001001010",
      "0001001011000000000000000000000001010111111000111111101101010010001001010110000" when "0001001011",
      "0001001100000000000000000000000001011010001111111111101101000010001110111010011" when "0001001100",
      "0001001101000000000000000000000001011100101000111111101100110010010100101000001" when "0001001101",
      "0001001110000000000000000000000001011111000011111111101100100010011010011111100" when "0001001110",
      "0001001111000000000000000000000001100001100000111111101100010010100000100000101" when "0001001111",
      "0001010000000000000000000000000001100011111111111111101100000010100110101011101" when "0001010000",
      "0001010001000000000000000000000001100110100000111111101011110010101101000000101" when "0001010001",
      "0001010010000000000000000000000001101001000011111111101011100010110011011111111" when "0001010010",
      "0001010011000000000000000000000001101011101000111111101011010010111010001001010" when "0001010011",
      "0001010100000000000000000000000001101110001111111111101011000011000000111101000" when "0001010100",
      "0001010101000000000000000000000001110000111000111111101010110011000111111011010" when "0001010101",
      "0001010110000000000000000000000001110011100011111111101010100011001111000100001" when "0001010110",
      "0001010111000000000000000000000001110110010000111111101010010011010110010111110" when "0001010111",
      "0001011000000000000000000000000001111000111111111111101010000011011101110110010" when "0001011000",
      "0001011001000000000000000000000001111011110000111111101001110011100101011111111" when "0001011001",
      "0001011010000000000000000000000001111110100011111111101001100011101101010100100" when "0001011010",
      "0001011011000000000000000000000010000001011000111111101001010011110101010100011" when "0001011011",
      "0001011100000000000000000000000010000100001111111111101001000011111101011111101" when "0001011100",
      "0001011101000000000000000000000010000111001000111111101000110100000101110110011" when "0001011101",
      "0001011110000000000000000000000010001010000011111111101000100100001110011000110" when "0001011110",
      "0001011111000000000000000000000010001101000000111111101000010100010111000111000" when "0001011111",
      "0001100000000000000000000000000010001111111111111111101000000100100000000001000" when "0001100000",
      "0001100001000000000000000000000010010011000000111111100111110100101001000111000" when "0001100001",
      "0001100010000000000000000000000010010110000011111111100111100100110010011001001" when "0001100010",
      "0001100011000000000000000000000010011001001000111111100111010100111011110111100" when "0001100011",
      "0001100100000000000000000000000010011100001111111111100111000101000101100010010" when "0001100100",
      "0001100101000000000000000000000010011111011000111111100110110101001111011001101" when "0001100101",
      "0001100110000000000000000000000010100010100011111111100110100101011001011101100" when "0001100110",
      "0001100111000000000000000000000010100101110000111111100110010101100011101110001" when "0001100111",
      "0001101000000000000000000000000010101000111111111111100110000101101110001011101" when "0001101000",
      "0001101001000000000000000000000010101100010000111111100101110101111000110110001" when "0001101001",
      "0001101010000000000000000000000010101111100011111111100101100110000011101101110" when "0001101010",
      "0001101011000000000000000000000010110010111000111111100101010110001110110010110" when "0001101011",
      "0001101100000000000000000000000010110110001111111111100101000110011010000101000" when "0001101100",
      "0001101101000000000000000000000010111001101000111111100100110110100101100100110" when "0001101101",
      "0001101110000000000000000000000010111101000011111111100100100110110001010010001" when "0001101110",
      "0001101111000000000000000000000011000000100000111111100100010110111101001101010" when "0001101111",
      "0001110000000000000000000000000011000011111111111111100100000111001001010110010" when "0001110000",
      "0001110001000000000000000000000011000111100000111111100011110111010101101101011" when "0001110001",
      "0001110010000000000000000000000011001011000011111111100011100111100010010010100" when "0001110010",
      "0001110011000000000000000000000011001110101000111111100011010111101111000101111" when "0001110011",
      "0001110100000000000000000000000011010010001111111111100011000111111100000111101" when "0001110100",
      "0001110101000000000000000000000011010101111000111111100010111000001001010111111" when "0001110101",
      "0001110110000000000000000000000011011001100011111111100010101000010110110110110" when "0001110110",
      "0001110111000000000000000000000011011101010000111111100010011000100100100100100" when "0001110111",
      "0001111000000000000000000000000011100000111111111111100010001000110010100001000" when "0001111000",
      "0001111001000000000000000000000011100100110000111111100001111001000000101100100" when "0001111001",
      "0001111010000000000000000000000011101000100011111111100001101001001111000111001" when "0001111010",
      "0001111011000000000000000000000011101100011000111111100001011001011101110001000" when "0001111011",
      "0001111100000000000000000000000011110000001111111111100001001001101100101010010" when "0001111100",
      "0001111101000000000000000000000011110100001000111111100000111001111011110011001" when "0001111101",
      "0001111110000000000000000000000011111000000011111111100000101010001011001011100" when "0001111110",
      "0001111111000000000000000000000011111100000000111111100000011010011010110011101" when "0001111111",
      "0010000000000000000000000000000011111111111111111111100000001010101010101011101" when "0010000000",
      "0010000001000000000000000000000100000100000000111111011111111010111010110011101" when "0010000001",
      "0010000010000000000000000000000100001000000011111111011111101011001011001011110" when "0010000010",
      "0010000011000000000000000000000100001100001000111111011111011011011011110100010" when "0010000011",
      "0010000100000000000000000000000100010000001111111111011111001011101100101101000" when "0010000100",
      "0010000101000000000000000000000100010100011000111111011110111011111101110110010" when "0010000101",
      "0010000110000000000000000000000100011000100011111111011110101100001111010000001" when "0010000110",
      "0010000111000000000000000000000100011100110000111111011110011100100000111010110" when "0010000111",
      "0010001000000000000000000000000100100000111111111111011110001100110010110110010" when "0010001000",
      "0010001001000000000000000000000100100101010000111111011101111101000101000010110" when "0010001001",
      "0010001010000000000000000000000100101001100011111111011101101101010111100000100" when "0010001010",
      "0010001011000000000000000000000100101101111000111111011101011101101010001111011" when "0010001011",
      "0010001100000000000000000000000100110010001111111111011101001101111101001111101" when "0010001100",
      "0010001101000000000000000000000100110110101000111111011100111110010000100001011" when "0010001101",
      "0010001110000000000000000000000100111011000011111111011100101110100100000100110" when "0010001110",
      "0010001111000000000000000000000100111111100000111111011100011110110111111010000" when "0010001111",
      "0010010000000000000000000000000101000011111111111111011100001111001100000001000" when "0010010000",
      "0010010001000000000000000000000101001000100000111111011011111111100000011010000" when "0010010001",
      "0010010010000000000000000000000101001101000011111111011011101111110101000101001" when "0010010010",
      "0010010011000000000000000000000101010001101000111111011011100000001010000010100" when "0010010011",
      "0010010100000000000000000000000101010110001111111111011011010000011111010010010" when "0010010100",
      "0010010101000000000000000000000101011010111000111111011011000000110100110100100" when "0010010101",
      "0010010110000000000000000000000101011111100011111111011010110001001010101001100" when "0010010110",
      "0010010111000000000000000000000101100100010000111111011010100001100000110001001" when "0010010111",
      "0010011000000000000000000000000101101000111111111111011010010001110111001011101" when "0010011000",
      "0010011001000000000000000000000101101101110000111111011010000010001101111001001" when "0010011001",
      "0010011010000000000000000000000101110010100011111111011001110010100100111001110" when "0010011010",
      "0010011011000000000000000000000101110111011000111111011001100010111100001101110" when "0010011011",
      "0010011100000000000000000000000101111100001111111111011001010011010011110101000" when "0010011100",
      "0010011101000000000000000000000110000001001000111111011001000011101011101111110" when "0010011101",
      "0010011110000000000000000000000110000110000011111111011000110100000011111110001" when "0010011110",
      "0010011111000000000000000000000110001011000000111111011000100100011100100000010" when "0010011111",
      "0010100000000000000000000000000110001111111111111111011000010100110101010110010" when "0010100000",
      "0010100001000000000000000000000110010101000000111111011000000101001110100000010" when "0010100001",
      "0010100010000000000000000000000110011010000011111111010111110101100111111110100" when "0010100010",
      "0010100011000000000000000000000110011111001000111111010111100110000001110000111" when "0010100011",
      "0010100100000000000000000000000110100100001111111111010111010110011011110111101" when "0010100100",
      "0010100101000000000000000000000110101001011000111111010111000110110110010010111" when "0010100101",
      "0010100110000000000000000000000110101110100011111111010110110111010001000010110" when "0010100110",
      "0010100111000000000000000000000110110011110000111111010110100111101100000111100" when "0010100111",
      "0010101000000000000000000000000110111000111111111111010110011000000111100001000" when "0010101000",
      "0010101001000000000000000000000110111110010000111111010110001000100011001111100" when "0010101001",
      "0010101010000000000000000000000111000011100011111111010101111000111111010011001" when "0010101010",
      "0010101011000000000000000000000111001000111000111111010101101001011011101100000" when "0010101011",
      "0010101100000000000000000000000111001110001111111111010101011001111000011010010" when "0010101100",
      "0010101101000000000000000000000111010011101000111111010101001010010101011110000" when "0010101101",
      "0010101110000000000000000000000111011001000011111111010100111010110010110111100" when "0010101110",
      "0010101111000000000000000000000111011110100000111111010100101011010000100110101" when "0010101111",
      "0010110000000000000000000000000111100011111111111111010100011011101110101011101" when "0010110000",
      "0010110001000000000000000000000111101001100000111111010100001100001101000110101" when "0010110001",
      "0010110010000000000000000000000111101111000011111111010011111100101011110111110" when "0010110010",
      "0010110011000000000000000000000111110100101000111111010011101101001010111111001" when "0010110011",
      "0010110100000000000000000000000111111010001111111111010011011101101010011101000" when "0010110100",
      "0010110101000000000000000000000111111111111000111111010011001110001010010001010" when "0010110101",
      "0010110110000000000000000000001000000101100011111111010010111110101010011100001" when "0010110110",
      "0010110111000000000000000000001000001011010000111111010010101111001010111101110" when "0010110111",
      "0010111000000000000000000000001000010000111111111111010010011111101011110110010" when "0010111000",
      "0010111001000000000000000000001000010110110000111111010010010000001101000101110" when "0010111001",
      "0010111010000000000000000000001000011100100011111111010010000000101110101100100" when "0010111010",
      "0010111011000000000000000000001000100010011000111111010001110001010000101010011" when "0010111011",
      "0010111100000000000000000000001000101000001111111111010001100001110010111111101" when "0010111100",
      "0010111101000000000000000000001000101110001000111111010001010010010101101100011" when "0010111101",
      "0010111110000000000000000000001000110100000011111111010001000010111000110000110" when "0010111110",
      "0010111111000000000000000000001000111010000000111111010000110011011100001100111" when "0010111111",
      "0011000000000000000000000000001000111111111111111111010000100100000000000001000" when "0011000000",
      "0011000001000000000000000000001001000110000000111111010000010100100100001101000" when "0011000001",
      "0011000010000000000000000000001001001100000011111111010000000101001000110001001" when "0011000010",
      "0011000011000000000000000000001001010010001000111111001111110101101101101101100" when "0011000011",
      "0011000100000000000000000000001001011000001111111111001111100110010011000010010" when "0011000100",
      "0011000101000000000000000000001001011110011000111111001111010110111000101111100" when "0011000101",
      "0011000110000000000000000000001001100100100011111111001111000111011110110101100" when "0011000110",
      "0011000111000000000000000000001001101010110000111111001110111000000101010100000" when "0011000111",
      "0011001000000000000000000000001001110000111111111111001110101000101100001011101" when "0011001000",
      "0011001001000000000000000000001001110111010000111111001110011001010011011100001" when "0011001001",
      "0011001010000000000000000000001001111101100011111111001110001001111011000101110" when "0011001010",
      "0011001011000000000000000000001010000011111000111111001101111010100011001000101" when "0011001011",
      "0011001100000000000000000000001010001010001111111111001101101011001011100100111" when "0011001100",
      "0011001101000000000000000000001010010000101000111111001101011011110100011010110" when "0011001101",
      "0011001110000000000000000000001010010111000011111111001101001100011101101010001" when "0011001110",
      "0011001111000000000000000000001010011101100000111111001100111101000111010011010" when "0011001111",
      "0011010000000000000000000000001010100011111111111111001100101101110001010110010" when "0011010000",
      "0011010001000000000000000000001010101010100000111111001100011110011011110011010" when "0011010001",
      "0011010010000000000000000000001010110001000011111111001100001111000110101010011" when "0011010010",
      "0011010011000000000000000000001010110111101000111111001011111111110001111011110" when "0011010011",
      "0011010100000000000000000000001010111110001111111111001011110000011101100111101" when "0011010100",
      "0011010101000000000000000000001011000100111000111111001011100001001001101101111" when "0011010101",
      "0011010110000000000000000000001011001011100011111111001011010001110110001110110" when "0011010110",
      "0011010111000000000000000000001011010010010000111111001011000010100011001010011" when "0011010111",
      "0011011000000000000000000000001011011000111111111111001010110011010000100000111" when "0011011000",
      "0011011001000000000000000000001011011111110000111111001010100011111110010010100" when "0011011001",
      "0011011010000000000000000000001011100110100011111111001010010100101100011111000" when "0011011010",
      "0011011011000000000000000000001011101101011000111111001010000101011011000111000" when "0011011011",
      "0011011100000000000000000000001011110100001111111111001001110110001010001010010" when "0011011100",
      "0011011101000000000000000000001011111011001000111111001001100110111001101001000" when "0011011101",
      "0011011110000000000000000000001100000010000011111111001001010111101001100011011" when "0011011110",
      "0011011111000000000000000000001100001001000000111111001001001000011001111001100" when "0011011111",
      "0011100000000000000000000000001100001111111111111111001000111001001010101011100" when "0011100000",
      "0011100001000000000000000000001100010111000000111111001000101001111011111001101" when "0011100001",
      "0011100010000000000000000000001100011110000011111111001000011010101101100011110" when "0011100010",
      "0011100011000000000000000000001100100101001000111111001000001011011111101010001" when "0011100011",
      "0011100100000000000000000000001100101100001111111111000111111100010010001100111" when "0011100100",
      "0011100101000000000000000000001100110011011000111111000111101101000101001100010" when "0011100101",
      "0011100110000000000000000000001100111010100011111111000111011101111000101000000" when "0011100110",
      "0011100111000000000000000000001101000001110000111111000111001110101100100000110" when "0011100111",
      "0011101000000000000000000000001101001000111111111111000110111111100000110110010" when "0011101000",
      "0011101001000000000000000000001101010000010000111111000110110000010101101000110" when "0011101001",
      "0011101010000000000000000000001101010111100011111111000110100001001010111000011" when "0011101010",
      "0011101011000000000000000000001101011110111000111111000110010010000000100101010" when "0011101011",
      "0011101100000000000000000000001101100110001111111111000110000010110110101111100" when "0011101100",
      "0011101101000000000000000000001101101101101000111111000101110011101101010111011" when "0011101101",
      "0011101110000000000000000000001101110101000011111111000101100100100100011100110" when "0011101110",
      "0011101111000000000000000000001101111100100000111111000101010101011011111111111" when "0011101111",
      "0011110000000000000000000000001110000011111111111111000101000110010100000000111" when "0011110000",
      "0011110001000000000000000000001110001011100000111111000100110111001100011111111" when "0011110001",
      "0011110010000000000000000000001110010011000011111111000100101000000101011101000" when "0011110010",
      "0011110011000000000000000000001110011010101000111111000100011000111110111000100" when "0011110011",
      "0011110100000000000000000000001110100010001111111111000100001001111000110010010" when "0011110100",
      "0011110101000000000000000000001110101001111000111111000011111010110011001010100" when "0011110101",
      "0011110110000000000000000000001110110001100011111111000011101011101110000001011" when "0011110110",
      "0011110111000000000000000000001110111001010000111111000011011100101001010111000" when "0011110111",
      "0011111000000000000000000000001111000000111111111111000011001101100101001011100" when "0011111000",
      "0011111001000000000000000000001111001000110000111111000010111110100001011111000" when "0011111001",
      "0011111010000000000000000000001111010000100011111111000010101111011110010001110" when "0011111010",
      "0011111011000000000000000000001111011000011000111111000010100000011011100011101" when "0011111011",
      "0011111100000000000000000000001111100000001111111111000010010001011001010100111" when "0011111100",
      "0011111101000000000000000000001111101000001000111111000010000010010111100101101" when "0011111101",
      "0011111110000000000000000000001111110000000011111111000001110011010110010110000" when "0011111110",
      "0011111111000000000000000000001111111000000000111111000001100100010101100110010" when "0011111111",
      "0100000000000000000000000000001111111111111111111111000001010101010101010110010" when "0100000000",
      "0100000001000000000000000000010000001000000000111111000001000110010101100110010" when "0100000001",
      "0100000010000000000000000000010000010000000011111111000000110111010110010110011" when "0100000010",
      "0100000011000000000000000000010000011000001000111111000000101000010111100110110" when "0100000011",
      "0100000100000000000000000000010000100000001111111111000000011001011001010111100" when "0100000100",
      "0100000101000000000000000000010000101000011000111111000000001010011011101000110" when "0100000101",
      "0100000110000000000000000000010000110000100011111110111111111011011110011010110" when "0100000110",
      "0100000111000000000000000000010000111000110000111110111111101100100001101101011" when "0100000111",
      "0100001000000000000000000000010001000000111111111110111111011101100101100000111" when "0100001000",
      "0100001001000000000000000000010001001001010000111110111111001110101001110101011" when "0100001001",
      "0100001010000000000000000000010001010001100011111110111110111111101110101011000" when "0100001010",
      "0100001011000000000000000000010001011001111000111110111110110000110100000010000" when "0100001011",
      "0100001100000000000000000000010001100010001111111110111110100001111001111010010" when "0100001100",
      "0100001101000000000000000000010001101010101000111110111110010011000000010100000" when "0100001101",
      "0100001110000000000000000000010001110011000011111110111110000100000111001111011" when "0100001110",
      "0100001111000000000000000000010001111011100000111110111101110101001110101100100" when "0100001111",
      "0100010000000000000000000000010010000011111111111110111101100110010110101011100" when "0100010000",
      "0100010001000000000000000000010010001100100000111110111101010111011111001100100" when "0100010001",
      "0100010010000000000000000000010010010101000011111110111101001000101000001111110" when "0100010010",
      "0100010011000000000000000000010010011101101000111110111100111001110001110101000" when "0100010011",
      "0100010100000000000000000000010010100110001111111110111100101010111011111100111" when "0100010100",
      "0100010101000000000000000000010010101110111000111110111100011100000110100111001" when "0100010101",
      "0100010110000000000000000000010010110111100011111110111100001101010001110100000" when "0100010110",
      "0100010111000000000000000000010011000000010000111110111011111110011101100011110" when "0100010111",
      "0100011000000000000000000000010011001000111111111110111011101111101001110110010" when "0100011000",
      "0100011001000000000000000000010011010001110000111110111011100000110110101011110" when "0100011001",
      "0100011010000000000000000000010011011010100011111110111011010010000100000100011" when "0100011010",
      "0100011011000000000000000000010011100011011000111110111011000011010010000000010" when "0100011011",
      "0100011100000000000000000000010011101100001111111110111010110100100000011111100" when "0100011100",
      "0100011101000000000000000000010011110101001000111110111010100101101111100010010" when "0100011101",
      "0100011110000000000000000000010011111110000011111110111010010110111111001000110" when "0100011110",
      "0100011111000000000000000000010100000111000000111110111010001000001111010010110" when "0100011111",
      "0100100000000000000000000000010100001111111111111110111001111001100000000000111" when "0100100000",
      "0100100001000000000000000000010100011001000000111110111001101010110001010010111" when "0100100001",
      "0100100010000000000000000000010100100010000011111110111001011100000011001001000" when "0100100010",
      "0100100011000000000000000000010100101011001000111110111001001101010101100011011" when "0100100011",
      "0100100100000000000000000000010100110100001111111110111000111110101000100010010" when "0100100100",
      "0100100101000000000000000000010100111101011000111110111000101111111100000101100" when "0100100101",
      "0100100110000000000000000000010101000110100011111110111000100001010000001101010" when "0100100110",
      "0100100111000000000000000000010101001111110000111110111000010010100100111010000" when "0100100111",
      "0100101000000000000000000000010101011000111111111110111000000011111010001011100" when "0100101000",
      "0100101001000000000000000000010101100010010000111110110111110101010000000010000" when "0100101001",
      "0100101010000000000000000000010101101011100011111110110111100110100110011101110" when "0100101010",
      "0100101011000000000000000000010101110100111000111110110111010111111101011110100" when "0100101011",
      "0100101100000000000000000000010101111110001111111110110111001001010101000100110" when "0100101100",
      "0100101101000000000000000000010110000111101000111110110110111010101101010000101" when "0100101101",
      "0100101110000000000000000000010110010001000011111110110110101100000110000010000" when "0100101110",
      "0100101111000000000000000000010110011010100000111110110110011101011111011001001" when "0100101111",
      "0100110000000000000000000000010110100011111111111110110110001110111001010110010" when "0100110000",
      "0100110001000000000000000000010110101101100000111110110110000000010011111001010" when "0100110001",
      "0100110010000000000000000000010110110111000011111110110101110001101111000010010" when "0100110010",
      "0100110011000000000000000000010111000000101000111110110101100011001010110001110" when "0100110011",
      "0100110100000000000000000000010111001010001111111110110101010100100111000111100" when "0100110100",
      "0100110101000000000000000000010111010011111000111110110101000110000100000011110" when "0100110101",
      "0100110110000000000000000000010111011101100011111110110100110111100001100110101" when "0100110110",
      "0100110111000000000000000000010111100111010000111110110100101000111111110000010" when "0100110111",
      "0100111000000000000000000000010111110000111111111110110100011010011110100000110" when "0100111000",
      "0100111001000000000000000000010111111010110000111110110100001011111101111000010" when "0100111001",
      "0100111010000000000000000000011000000100100011111110110011111101011101110111000" when "0100111010",
      "0100111011000000000000000000011000001110011000111110110011101110111110011100111" when "0100111011",
      "0100111100000000000000000000011000011000001111111110110011100000011111101010001" when "0100111100",
      "0100111101000000000000000000011000100010001000111110110011010010000001011111000" when "0100111101",
      "0100111110000000000000000000011000101100000011111110110011000011100011111011010" when "0100111110",
      "0100111111000000000000000000011000110110000000111110110010110101000110111111100" when "0100111111",
      "0101000000000000000000000000011000111111111111111110110010100110101010101011100" when "0101000000",
      "0101000001000000000000000000011001001010000000111110110010011000001110111111100" when "0101000001",
      "0101000010000000000000000000011001010100000011111110110010001001110011111011101" when "0101000010",
      "0101000011000000000000000000011001011110001000111110110001111011011001100000000" when "0101000011",
      "0101000100000000000000000000011001101000001111111110110001101100111111101100110" when "0101000100",
      "0101000101000000000000000000011001110010011000111110110001011110100110100010000" when "0101000101",
      "0101000110000000000000000000011001111100100011111110110001010000001110000000000" when "0101000110",
      "0101000111000000000000000000011010000110110000111110110001000001110110000110101" when "0101000111",
      "0101001000000000000000000000011010010000111111111110110000110011011110110110001" when "0101001000",
      "0101001001000000000000000000011010011011010000111110110000100101001000001110101" when "0101001001",
      "0101001010000000000000000000011010100101100011111110110000010110110010010000010" when "0101001010",
      "0101001011000000000000000000011010101111111000111110110000001000011100111011010" when "0101001011",
      "0101001100000000000000000000011010111010001111111110101111111010001000001111100" when "0101001100",
      "0101001101000000000000000000011011000100101000111110101111101011110100001101010" when "0101001101",
      "0101001110000000000000000000011011001111000011111110101111011101100000110100101" when "0101001110",
      "0101001111000000000000000000011011011001100000111110101111001111001110000101110" when "0101001111",
      "0101010000000000000000000000011011100011111111111110101111000000111100000000110" when "0101010000",
      "0101010001000000000000000000011011101110100000111110101110110010101010100101110" when "0101010001",
      "0101010010000000000000000000011011111001000011111110101110100100011001110101000" when "0101010010",
      "0101010011000000000000000000011100000011101000111110101110010110001001101110011" when "0101010011",
      "0101010100000000000000000000011100001110001111111110101110000111111010010010001" when "0101010100",
      "0101010101000000000000000000011100011000111000111110101101111001101011100000011" when "0101010101",
      "0101010110000000000000000000011100100011100011111110101101101011011101011001010" when "0101010110",
      "0101010111000000000000000000011100101110010000111110101101011101001111111101000" when "0101010111",
      "0101011000000000000000000000011100111000111111111110101101001111000011001011100" when "0101011000",
      "0101011001000000000000000000011101000011110000111110101101000000110111000101000" when "0101011001",
      "0101011010000000000000000000011101001110100011111110101100110010101011101001101" when "0101011010",
      "0101011011000000000000000000011101011001011000111110101100100100100000111001100" when "0101011011",
      "0101011100000000000000000000011101100100001111111110101100010110010110110100110" when "0101011100",
      "0101011101000000000000000000011101101111001000111110101100001000001101011011100" when "0101011101",
      "0101011110000000000000000000011101111010000011111110101011111010000100101110000" when "0101011110",
      "0101011111000000000000000000011110000101000000111110101011101011111100101100000" when "0101011111",
      "0101100000000000000000000000011110001111111111111110101011011101110101010110001" when "0101100000",
      "0101100001000000000000000000011110011011000000111110101011001111101110101100001" when "0101100001",
      "0101100010000000000000000000011110100110000011111110101011000001101000101110010" when "0101100010",
      "0101100011000000000000000000011110110001001000111110101010110011100011011100110" when "0101100011",
      "0101100100000000000000000000011110111100001111111110101010100101011110110111100" when "0101100100",
      "0101100101000000000000000000011111000111011000111110101010010111011010111110110" when "0101100101",
      "0101100110000000000000000000011111010010100011111110101010001001010111110010101" when "0101100110",
      "0101100111000000000000000000011111011101110000111110101001111011010101010011010" when "0101100111",
      "0101101000000000000000000000011111101000111111111110101001101101010011100000110" when "0101101000",
      "0101101001000000000000000000011111110100010000111110101001011111010010011011010" when "0101101001",
      "0101101010000000000000000000011111111111100011111110101001010001010010000011000" when "0101101010",
      "0101101011000000000000000000100000001010111000111110101001000011010010010111110" when "0101101011",
      "0101101100000000000000000000100000010110001111111110101000110101010011011010000" when "0101101100",
      "0101101101000000000000000000100000100001101000111110101000100111010101001001111" when "0101101101",
      "0101101110000000000000000000100000101101000011111110101000011001010111100111010" when "0101101110",
      "0101101111000000000000000000100000111000100000111110101000001011011010110010011" when "0101101111",
      "0101110000000000000000000000100001000011111111111110100111111101011110101011100" when "0101110000",
      "0101110001000000000000000000100001001111100000111110100111101111100011010010100" when "0101110001",
      "0101110010000000000000000000100001011011000011111110100111100001101000100111100" when "0101110010",
      "0101110011000000000000000000100001100110101000111110100111010011101110101011000" when "0101110011",
      "0101110100000000000000000000100001110010001111111110100111000101110101011100110" when "0101110100",
      "0101110101000000000000000000100001111101111000111110100110110111111100111101000" when "0101110101",
      "0101110110000000000000000000100010001001100011111110100110101010000101001100000" when "0101110110",
      "0101110111000000000000000000100010010101010000111110100110011100001110001001100" when "0101110111",
      "0101111000000000000000000000100010100000111111111110100110001110010111110110000" when "0101111000",
      "0101111001000000000000000000100010101100110000111110100110000000100010010001100" when "0101111001",
      "0101111010000000000000000000100010111000100011111110100101110010101101011100010" when "0101111010",
      "0101111011000000000000000000100011000100011000111110100101100100111001010110001" when "0101111011",
      "0101111100000000000000000000100011010000001111111110100101010111000101111111011" when "0101111100",
      "0101111101000000000000000000100011011100001000111110100101001001010011011000010" when "0101111101",
      "0101111110000000000000000000100011101000000011111110100100111011100001100000100" when "0101111110",
      "0101111111000000000000000000100011110100000000111110100100101101110000011000110" when "0101111111",
      "0110000000000000000000000000100011111111111111111110100100100000000000000000110" when "0110000000",
      "0110000001000000000000000000100100001100000000111110100100010010010000011000110" when "0110000001",
      "0110000010000000000000000000100100011000000011111110100100000100100001100000111" when "0110000010",
      "0110000011000000000000000000100100100100001000111110100011110110110011011001010" when "0110000011",
      "0110000100000000000000000000100100110000001111111110100011101001000110000010000" when "0110000100",
      "0110000101000000000000000000100100111100011000111110100011011011011001011011010" when "0110000101",
      "0110000110000000000000000000100101001000100011111110100011001101101101100101010" when "0110000110",
      "0110000111000000000000000000100101010100110000111110100011000000000010011111111" when "0110000111",
      "0110001000000000000000000000100101100000111111111110100010110010011000001011011" when "0110001000",
      "0110001001000000000000000000100101101101010000111110100010100100101110100111111" when "0110001001",
      "0110001010000000000000000000100101111001100011111110100010010111000101110101100" when "0110001010",
      "0110001011000000000000000000100110000101111000111110100010001001011101110100100" when "0110001011",
      "0110001100000000000000000000100110010010001111111110100001111011110110100100110" when "0110001100",
      "0110001101000000000000000000100110011110101000111110100001101110010000000110100" when "0110001101",
      "0110001110000000000000000000100110101011000011111110100001100000101010011001111" when "0110001110",
      "0110001111000000000000000000100110110111100000111110100001010011000101011111000" when "0110001111",
      "0110010000000000000000000000100111000011111111111110100001000101100001010110000" when "0110010000",
      "0110010001000000000000000000100111010000100000111110100000110111111101111111000" when "0110010001",
      "0110010010000000000000000000100111011101000011111110100000101010011011011010010" when "0110010010",
      "0110010011000000000000000000100111101001101000111110100000011100111001100111101" when "0110010011",
      "0110010100000000000000000000100111110110001111111110100000001111011000100111011" when "0110010100",
      "0110010101000000000000000000101000000010111000111110100000000001111000011001101" when "0110010101",
      "0110010110000000000000000000101000001111100011111110011111110100011000111110100" when "0110010110",
      "0110010111000000000000000000101000011100010000111110011111100110111010010110010" when "0110010111",
      "0110011000000000000000000000101000101000111111111110011111011001011100100000110" when "0110011000",
      "0110011001000000000000000000101000110101110000111110011111001011111111011110010" when "0110011001",
      "0110011010000000000000000000101001000010100011111110011110111110100011001110111" when "0110011010",
      "0110011011000000000000000000101001001111011000111110011110110001000111110010110" when "0110011011",
      "0110011100000000000000000000101001011100001111111110011110100011101101001010000" when "0110011100",
      "0110011101000000000000000000101001101001001000111110011110010110010011010100110" when "0110011101",
      "0110011110000000000000000000101001110110000011111110011110001000111010010011010" when "0110011110",
      "0110011111000000000000000000101010000011000000111110011101111011100010000101010" when "0110011111",
      "0110100000000000000000000000101010001111111111111110011101101110001010101011011" when "0110100000",
      "0110100001000000000000000000101010011101000000111110011101100000110100000101011" when "0110100001",
      "0110100010000000000000000000101010101010000011111110011101010011011110010011100" when "0110100010",
      "0110100011000000000000000000101010110111001000111110011101000110001001010110000" when "0110100011",
      "0110100100000000000000000000101011000100001111111110011100111000110101001100110" when "0110100100",
      "0110100101000000000000000000101011010001011000111110011100101011100001111000000" when "0110100101",
      "0110100110000000000000000000101011011110100011111110011100011110001111010111110" when "0110100110",
      "0110100111000000000000000000101011101011110000111110011100010000111101101100100" when "0110100111",
      "0110101000000000000000000000101011111000111111111110011100000011101100110110000" when "0110101000",
      "0110101001000000000000000000101100000110010000111110011011110110011100110100100" when "0110101001",
      "0110101010000000000000000000101100010011100011111110011011101001001101101000010" when "0110101010",
      "0110101011000000000000000000101100100000111000111110011011011011111111010001000" when "0110101011",
      "0110101100000000000000000000101100101110001111111110011011001110110001101111010" when "0110101100",
      "0110101101000000000000000000101100111011101000111110011011000001100101000011001" when "0110101101",
      "0110101110000000000000000000101101001001000011111110011010110100011001001100100" when "0110101110",
      "0110101111000000000000000000101101010110100000111110011010100111001110001011101" when "0110101111",
      "0110110000000000000000000000101101100011111111111110011010011010000100000000110" when "0110110000",
      "0110110001000000000000000000101101110001100000111110011010001100111010101011110" when "0110110001",
      "0110110010000000000000000000101101111111000011111110011001111111110010001100110" when "0110110010",
      "0110110011000000000000000000101110001100101000111110011001110010101010100100010" when "0110110011",
      "0110110100000000000000000000101110011010001111111110011001100101100011110010000" when "0110110100",
      "0110110101000000000000000000101110100111111000111110011001011000011101110110010" when "0110110101",
      "0110110110000000000000000000101110110101100011111110011001001011011000110001001" when "0110110110",
      "0110110111000000000000000000101111000011010000111110011000111110010100100010110" when "0110110111",
      "0110111000000000000000000000101111010000111111111110011000110001010001001011010" when "0110111000",
      "0110111001000000000000000000101111011110110000111110011000100100001110101010110" when "0110111001",
      "0110111010000000000000000000101111101100100011111110011000010111001101000001100" when "0110111010",
      "0110111011000000000000000000101111111010011000111110011000001010001100001111011" when "0110111011",
      "0110111100000000000000000000110000001000001111111110010111111101001100010100101" when "0110111100",
      "0110111101000000000000000000110000010110001000111110010111110000001101010001100" when "0110111101",
      "0110111110000000000000000000110000100100000011111110010111100011001111000101110" when "0110111110",
      "0110111111000000000000000000110000110010000000111110010111010110010001110010000" when "0110111111",
      "0111000000000000000000000000110000111111111111111110010111001001010101010110000" when "0111000000",
      "0111000001000000000000000000110001001110000000111110010110111100011001110010000" when "0111000001",
      "0111000010000000000000000000110001011100000011111110010110101111011111000110001" when "0111000010",
      "0111000011000000000000000000110001101010001000111110010110100010100101010010100" when "0111000011",
      "0111000100000000000000000000110001111000001111111110010110010101101100010111010" when "0111000100",
      "0111000101000000000000000000110010000110011000111110010110001000110100010100100" when "0111000101",
      "0111000110000000000000000000110010010100100011111110010101111011111101001010100" when "0111000110",
      "0111000111000000000000000000110010100010110000111110010101101111000110111001001" when "0111000111",
      "0111001000000000000000000000110010110000111111111110010101100010010001100000101" when "0111001000",
      "0111001001000000000000000000110010111111010000111110010101010101011101000001001" when "0111001001",
      "0111001010000000000000000000110011001101100011111110010101001000101001011010110" when "0111001010",
      "0111001011000000000000000000110011011011111000111110010100111011110110101101110" when "0111001011",
      "0111001100000000000000000000110011101010001111111110010100101111000100111010000" when "0111001100",
      "0111001101000000000000000000110011111000101000111110010100100010010011111111110" when "0111001101",
      "0111001110000000000000000000110100000111000011111110010100010101100011111111001" when "0111001110",
      "0111001111000000000000000000110100010101100000111110010100001000110100111000010" when "0111001111",
      "0111010000000000000000000000110100100011111111111110010011111100000110101011010" when "0111010000",
      "0111010001000000000000000000110100110010100000111110010011101111011001011000010" when "0111010001",
      "0111010010000000000000000000110101000001000011111110010011100010101100111111100" when "0111010010",
      "0111010011000000000000000000110101001111101000111110010011010110000001100000110" when "0111010011",
      "0111010100000000000000000000110101011110001111111110010011001001010110111100101" when "0111010100",
      "0111010101000000000000000000110101101100111000111110010010111100101101010010111" when "0111010101",
      "0111010110000000000000000000110101111011100011111110010010110000000100100011110" when "0111010110",
      "0111010111000000000000000000110110001010010000111110010010100011011100101111100" when "0111010111",
      "0111011000000000000000000000110110011000111111111110010010010110110101110110000" when "0111011000",
      "0111011001000000000000000000110110100111110000111110010010001010001111110111100" when "0111011001",
      "0111011010000000000000000000110110110110100011111110010001111101101010110100001" when "0111011010",
      "0111011011000000000000000000110111000101011000111110010001110001000110101100000" when "0111011011",
      "0111011100000000000000000000110111010100001111111110010001100100100011011111010" when "0111011100",
      "0111011101000000000000000000110111100011001000111110010001011000000001001110000" when "0111011101",
      "0111011110000000000000000000110111110010000011111110010001001011011111111000100" when "0111011110",
      "0111011111000000000000000000111000000001000000111110010000111110111111011110100" when "0111011111",
      "0111100000000000000000000000111000001111111111111110010000110010100000000000100" when "0111100000",
      "0111100001000000000000000000111000011111000000111110010000100110000001011110101" when "0111100001",
      "0111100010000000000000000000111000101110000011111110010000011001100011111000110" when "0111100010",
      "0111100011000000000000000000111000111101001000111110010000001101000111001111001" when "0111100011",
      "0111100100000000000000000000111001001100001111111110010000000000101011100010000" when "0111100100",
      "0111100101000000000000000000111001011011011000111110001111110100010000110001010" when "0111100101",
      "0111100110000000000000000000111001101010100011111110001111100111110110111101000" when "0111100110",
      "0111100111000000000000000000111001111001110000111110001111011011011110000101110" when "0111100111",
      "0111101000000000000000000000111010001000111111111110001111001111000110001011010" when "0111101000",
      "0111101001000000000000000000111010011000010000111110001111000010101111001101110" when "0111101001",
      "0111101010000000000000000000111010100111100011111110001110110110011001001101011" when "0111101010",
      "0111101011000000000000000000111010110110111000111110001110101010000100001010010" when "0111101011",
      "0111101100000000000000000000111011000110001111111110001110011101110000000100100" when "0111101100",
      "0111101101000000000000000000111011010101101000111110001110010001011100111100010" when "0111101101",
      "0111101110000000000000000000111011100101000011111110001110000101001010110001110" when "0111101110",
      "0111101111000000000000000000111011110100100000111110001101111000111001100100111" when "0111101111",
      "0111110000000000000000000000111100000011111111111110001101101100101001010101111" when "0111110000",
      "0111110001000000000000000000111100010011100000111110001101100000011010000101000" when "0111110001",
      "0111110010000000000000000000111100100011000011111110001101010100001011110010000" when "0111110010",
      "0111110011000000000000000000111100110010101000111110001101000111111110011101100" when "0111110011",
      "0111110100000000000000000000111101000010001111111110001100111011110010000111010" when "0111110100",
      "0111110101000000000000000000111101010001111000111110001100101111100110101111100" when "0111110101",
      "0111110110000000000000000000111101100001100011111110001100100011011100010110011" when "0111110110",
      "0111110111000000000000000000111101110001010000111110001100010111010010111100000" when "0111110111",
      "0111111000000000000000000000111110000000111111111110001100001011001010100000100" when "0111111000",
      "0111111001000000000000000000111110010000110000111110001011111111000011000100000" when "0111111001",
      "0111111010000000000000000000111110100000100011111110001011110010111100100110110" when "0111111010",
      "0111111011000000000000000000111110110000011000111110001011100110110111001000101" when "0111111011",
      "0111111100000000000000000000111111000000001111111110001011011010110010101001111" when "0111111100",
      "0111111101000000000000000000111111010000001000111110001011001110101111001010101" when "0111111101",
      "0111111110000000000000000000111111100000000011111110001011000010101100101011000" when "0111111110",
      "0111111111000000000000000000111111110000000000111110001010110110101011001011010" when "0111111111",
      "1000000000000000000000000000111111111111111111111110001010101010101010101011010" when "1000000000",
      "1000000001000000000000000001000000010000000000111110001010011110101011001011010" when "1000000001",
      "1000000010000000000000000001000000100000000011111110001010010010101100101011011" when "1000000010",
      "1000000011000000000000000001000000110000001000111110001010000110101111001011110" when "1000000011",
      "1000000100000000000000000001000001000000001111111110001001111010110010101100100" when "1000000100",
      "1000000101000000000000000001000001010000011000111110001001101110110111001101110" when "1000000101",
      "1000000110000000000000000001000001100000100011111110001001100010111100101111110" when "1000000110",
      "1000000111000000000000000001000001110000110000111110001001010111000011010010011" when "1000000111",
      "1000001000000000000000000001000010000000111111111110001001001011001010110101111" when "1000001000",
      "1000001001000000000000000001000010010001010000111110001000111111010011011010011" when "1000001001",
      "1000001010000000000000000001000010100001100011111110001000110011011101000000000" when "1000001010",
      "1000001011000000000000000001000010110001111000111110001000100111100111100110111" when "1000001011",
      "1000001100000000000000000001000011000010001111111110001000011011110011001111001" when "1000001100",
      "1000001101000000000000000001000011010010101000111110001000001111111111111001000" when "1000001101",
      "1000001110000000000000000001000011100011000011111110001000000100001101100100011" when "1000001110",
      "1000001111000000000000000001000011110011100000111110000111111000011100010001100" when "1000001111",
      "1000010000000000000000000001000100000011111111111110000111101100101100000000100" when "1000010000",
      "1000010001000000000000000001000100010100100000111110000111100000111100110001100" when "1000010001",
      "1000010010000000000000000001000100100101000011111110000111010101001110100100101" when "1000010010",
      "1000010011000000000000000001000100110101101000111110000111001001100001011010000" when "1000010011",
      "1000010100000000000000000001000101000110001111111110000110111101110101010001111" when "1000010100",
      "1000010101000000000000000001000101010110111000111110000110110010001010001100001" when "1000010101",
      "1000010110000000000000000001000101100111100011111110000110100110100000001001000" when "1000010110",
      "1000010111000000000000000001000101111000010000111110000110011010110111001000101" when "1000010111",
      "1000011000000000000000000001000110001000111111111110000110001111001111001011001" when "1000011000",
      "1000011001000000000000000001000110011001110000111110000110000011101000010000101" when "1000011001",
      "1000011010000000000000000001000110101010100011111110000101111000000010011001011" when "1000011010",
      "1000011011000000000000000001000110111011011000111110000101101100011101100101010" when "1000011011",
      "1000011100000000000000000001000111001100001111111110000101100000111001110100100" when "1000011100",
      "1000011101000000000000000001000111011101001000111110000101010101010111000111010" when "1000011101",
      "1000011110000000000000000001000111101110000011111110000101001001110101011101101" when "1000011110",
      "1000011111000000000000000001000111111111000000111110000100111110010100110111110" when "1000011111",
      "1000100000000000000000000001001000001111111111111110000100110010110101010101110" when "1000100000",
      "1000100001000000000000000001001000100001000000111110000100100111010110110111111" when "1000100001",
      "1000100010000000000000000001001000110010000011111110000100011011111001011110000" when "1000100010",
      "1000100011000000000000000001001001000011001000111110000100010000011101001000011" when "1000100011",
      "1000100100000000000000000001001001010100001111111110000100000101000001110111001" when "1000100100",
      "1000100101000000000000000001001001100101011000111110000011111001100111101010011" when "1000100101",
      "1000100110000000000000000001001001110110100011111110000011101110001110100010010" when "1000100110",
      "1000100111000000000000000001001010000111110000111110000011100010110110011111000" when "1000100111",
      "1000101000000000000000000001001010011000111111111110000011010111011111100000100" when "1000101000",
      "1000101001000000000000000001001010101010010000111110000011001100001001100111000" when "1000101001",
      "1000101010000000000000000001001010111011100011111110000011000000110100110010101" when "1000101010",
      "1000101011000000000000000001001011001100111000111110000010110101100001000011100" when "1000101011",
      "1000101100000000000000000001001011011110001111111110000010101010001110011001110" when "1000101100",
      "1000101101000000000000000001001011101111101000111110000010011110111100110101100" when "1000101101",
      "1000101110000000000000000001001100000001000011111110000010010011101100010111000" when "1000101110",
      "1000101111000000000000000001001100010010100000111110000010001000011100111110001" when "1000101111",
      "1000110000000000000000000001001100100011111111111110000001111101001110101011001" when "1000110000",
      "1000110001000000000000000001001100110101100000111110000001110010000001011110001" when "1000110001",
      "1000110010000000000000000001001101000111000011111110000001100110110101010111010" when "1000110010",
      "1000110011000000000000000001001101011000101000111110000001011011101010010110101" when "1000110011",
      "1000110100000000000000000001001101101010001111111110000001010000100000011100100" when "1000110100",
      "1000110101000000000000000001001101111011111000111110000001000101010111101000110" when "1000110101",
      "1000110110000000000000000001001110001101100011111110000000111010001111111011101" when "1000110110",
      "1000110111000000000000000001001110011111010000111110000000101111001001010101010" when "1000110111",
      "1000111000000000000000000001001110110000111111111110000000100100000011110101110" when "1000111000",
      "1000111001000000000000000001001111000010110000111110000000011000111111011101010" when "1000111001",
      "1000111010000000000000000001001111010100100011111110000000001101111100001011111" when "1000111010",
      "1000111011000000000000000001001111100110011000111110000000000010111010000001111" when "1000111011",
      "1000111100000000000000000001001111111000001111111101111111110111111000111111001" when "1000111100",
      "1000111101000000000000000001010000001010001000111101111111101100111001000011111" when "1000111101",
      "1000111110000000000000000001010000011100000011111101111111100001111010010000010" when "1000111110",
      "1000111111000000000000000001010000101110000000111101111111010110111100100100011" when "1000111111",
      "1001000000000000000000000001010000111111111111111101111111001100000000000000011" when "1001000000",
      "1001000001000000000000000001010001010010000000111101111111000001000100100100011" when "1001000001",
      "1001000010000000000000000001010001100100000011111101111110110110001010010000101" when "1001000010",
      "1001000011000000000000000001010001110110001000111101111110101011010001000101000" when "1001000011",
      "1001000100000000000000000001010010001000001111111101111110100000011001000001110" when "1001000100",
      "1001000101000000000000000001010010011010011000111101111110010101100010000111000" when "1001000101",
      "1001000110000000000000000001010010101100100011111101111110001010101100010100111" when "1001000110",
      "1001000111000000000000000001010010111110110000111101111101111111110111101011100" when "1001000111",
      "1001001000000000000000000001010011010000111111111101111101110101000100001011001" when "1001001000",
      "1001001001000000000000000001010011100011010000111101111101101010010001110011101" when "1001001001",
      "1001001010000000000000000001010011110101100011111101111101011111100000100101010" when "1001001010",
      "1001001011000000000000000001010100000111111000111101111101010100110000100000001" when "1001001011",
      "1001001100000000000000000001010100011010001111111101111101001010000001100100011" when "1001001100",
      "1001001101000000000000000001010100101100101000111101111100111111010011110010001" when "1001001101",
      "1001001110000000000000000001010100111111000011111101111100110100100111001001100" when "1001001110",
      "1001001111000000000000000001010101010001100000111101111100101001111011101010110" when "1001001111",
      "1001010000000000000000000001010101100011111111111101111100011111010001010101110" when "1001010000",
      "1001010001000000000000000001010101110110100000111101111100010100101000001010110" when "1001010001",
      "1001010010000000000000000001010110001001000011111101111100001010000000001001111" when "1001010010",
      "1001010011000000000000000001010110011011101000111101111011111111011001010011010" when "1001010011",
      "1001010100000000000000000001010110101110001111111101111011110100110011100111000" when "1001010100",
      "1001010101000000000000000001010111000000111000111101111011101010001111000101011" when "1001010101",
      "1001010110000000000000000001010111010011100011111101111011011111101011101110010" when "1001010110",
      "1001010111000000000000000001010111100110010000111101111011010101001001100001111" when "1001010111",
      "1001011000000000000000000001010111111000111111111101111011001010101000100000011" when "1001011000",
      "1001011001000000000000000001011000001011110000111101111011000000001000101001111" when "1001011001",
      "1001011010000000000000000001011000011110100011111101111010110101101001111110100" when "1001011010",
      "1001011011000000000000000001011000110001011000111101111010101011001100011110011" when "1001011011",
      "1001011100000000000000000001011001000100001111111101111010100000110000001001110" when "1001011100",
      "1001011101000000000000000001011001010111001000111101111010010110010101000000100" when "1001011101",
      "1001011110000000000000000001011001101010000011111101111010001011111011000010111" when "1001011110",
      "1001011111000000000000000001011001111101000000111101111010000001100010010001000" when "1001011111",
      "1001100000000000000000000001011010001111111111111101111001110111001010101011000" when "1001100000",
      "1001100001000000000000000001011010100011000000111101111001101100110100010001000" when "1001100001",
      "1001100010000000000000000001011010110110000011111101111001100010011111000011001" when "1001100010",
      "1001100011000000000000000001011011001001001000111101111001011000001011000001101" when "1001100011",
      "1001100100000000000000000001011011011100001111111101111001001101111000001100011" when "1001100100",
      "1001100101000000000000000001011011101111011000111101111001000011100110100011101" when "1001100101",
      "1001100110000000000000000001011100000010100011111101111000111001010110000111100" when "1001100110",
      "1001100111000000000000000001011100010101110000111101111000101111000110111000001" when "1001100111",
      "1001101000000000000000000001011100101000111111111101111000100100111000110101101" when "1001101000",
      "1001101001000000000000000001011100111100010000111101111000011010101100000000010" when "1001101001",
      "1001101010000000000000000001011101001111100011111101111000010000100000010111111" when "1001101010",
      "1001101011000000000000000001011101100010111000111101111000000110010101111100110" when "1001101011",
      "1001101100000000000000000001011101110110001111111101110111111100001100101111000" when "1001101100",
      "1001101101000000000000000001011110001001101000111101110111110010000100101110110" when "1001101101",
      "1001101110000000000000000001011110011101000011111101110111100111111101111100001" when "1001101110",
      "1001101111000000000000000001011110110000100000111101110111011101111000010111010" when "1001101111",
      "1001110000000000000000000001011111000011111111111101110111010011110100000000011" when "1001110000",
      "1001110001000000000000000001011111010111100000111101110111001001110000110111011" when "1001110001",
      "1001110010000000000000000001011111101011000011111101110110111111101110111100100" when "1001110010",
      "1001110011000000000000000001011111111110101000111101110110110101101110001111111" when "1001110011",
      "1001110100000000000000000001100000010010001111111101110110101011101110110001101" when "1001110100",
      "1001110101000000000000000001100000100101111000111101110110100001110000100001111" when "1001110101",
      "1001110110000000000000000001100000111001100011111101110110010111110011100000111" when "1001110110",
      "1001110111000000000000000001100001001101010000111101110110001101110111101110100" when "1001110111",
      "1001111000000000000000000001100001100000111111111101110110000011111101001011000" when "1001111000",
      "1001111001000000000000000001100001110100110000111101110101111010000011110110100" when "1001111001",
      "1001111010000000000000000001100010001000100011111101110101110000001011110001001" when "1001111010",
      "1001111011000000000000000001100010011100011000111101110101100110010100111011000" when "1001111011",
      "1001111100000000000000000001100010110000001111111101110101011100011111010100010" when "1001111100",
      "1001111101000000000000000001100011000100001000111101110101010010101010111101001" when "1001111101",
      "1001111110000000000000000001100011011000000011111101110101001000110111110101100" when "1001111110",
      "1001111111000000000000000001100011101100000000111101110100111111000101111101101" when "1001111111",
      "1010000000000000000000000001100011111111111111111101110100110101010101010101101" when "1010000000",
      "1010000001000000000000000001100100010100000000111101110100101011100101111101101" when "1010000001",
      "1010000010000000000000000001100100101000000011111101110100100001110111110101110" when "1010000010",
      "1010000011000000000000000001100100111100001000111101110100011000001010111110001" when "1010000011",
      "1010000100000000000000000001100101010000001111111101110100001110011111010111000" when "1010000100",
      "1010000101000000000000000001100101100100011000111101110100000100110101000000010" when "1010000101",
      "1010000110000000000000000001100101111000100011111101110011111011001011111010001" when "1010000110",
      "1010000111000000000000000001100110001100110000111101110011110001100100000100110" when "1010000111",
      "1010001000000000000000000001100110100000111111111101110011100111111101100000010" when "1010001000",
      "1010001001000000000000000001100110110101010000111101110011011110011000001100110" when "1010001001",
      "1010001010000000000000000001100111001001100011111101110011010100110100001010100" when "1010001010",
      "1010001011000000000000000001100111011101111000111101110011001011010001011001011" when "1010001011",
      "1010001100000000000000000001100111110010001111111101110011000001101111111001101" when "1010001100",
      "1010001101000000000000000001101000000110101000111101110010111000001111101011011" when "1010001101",
      "1010001110000000000000000001101000011011000011111101110010101110110000101110110" when "1010001110",
      "1010001111000000000000000001101000101111100000111101110010100101010011000011111" when "1010001111",
      "1010010000000000000000000001101001000011111111111101110010011011110110101010111" when "1010010000",
      "1010010001000000000000000001101001011000100000111101110010010010011011100100000" when "1010010001",
      "1010010010000000000000000001101001101101000011111101110010001001000001101111001" when "1010010010",
      "1010010011000000000000000001101010000001101000111101110001111111101001001100100" when "1010010011",
      "1010010100000000000000000001101010010110001111111101110001110110010001111100010" when "1010010100",
      "1010010101000000000000000001101010101010111000111101110001101100111011111110100" when "1010010101",
      "1010010110000000000000000001101010111111100011111101110001100011100111010011011" when "1010010110",
      "1010010111000000000000000001101011010100010000111101110001011010010011111011000" when "1010010111",
      "1010011000000000000000000001101011101000111111111101110001010001000001110101101" when "1010011000",
      "1010011001000000000000000001101011111101110000111101110001000111110001000011001" when "1010011001",
      "1010011010000000000000000001101100010010100011111101110000111110100001100011110" when "1010011010",
      "1010011011000000000000000001101100100111011000111101110000110101010011010111101" when "1010011011",
      "1010011100000000000000000001101100111100001111111101110000101100000110011110111" when "1010011100",
      "1010011101000000000000000001101101010001001000111101110000100010111010111001101" when "1010011101",
      "1010011110000000000000000001101101100110000011111101110000011001110000101000001" when "1010011110",
      "1010011111000000000000000001101101111011000000111101110000010000100111101010010" when "1010011111",
      "1010100000000000000000000001101110001111111111111101110000000111100000000000010" when "1010100000",
      "1010100001000000000000000001101110100101000000111101101111111110011001101010010" when "1010100001",
      "1010100010000000000000000001101110111010000011111101101111110101010100101000011" when "1010100010",
      "1010100011000000000000000001101111001111001000111101101111101100010000111010110" when "1010100011",
      "1010100100000000000000000001101111100100001111111101101111100011001110100001100" when "1010100100",
      "1010100101000000000000000001101111111001011000111101101111011010001101011100111" when "1010100101",
      "1010100110000000000000000001110000001110100011111101101111010001001101101100110" when "1010100110",
      "1010100111000000000000000001110000100011110000111101101111001000001111010001011" when "1010100111",
      "1010101000000000000000000001110000111000111111111101101110111111010010001010111" when "1010101000",
      "1010101001000000000000000001110001001110010000111101101110110110010110011001011" when "1010101001",
      "1010101010000000000000000001110001100011100011111101101110101101011011111101000" when "1010101010",
      "1010101011000000000000000001110001111000111000111101101110100100100010110110000" when "1010101011",
      "1010101100000000000000000001110010001110001111111101101110011011101011000100010" when "1010101100",
      "1010101101000000000000000001110010100011101000111101101110010010110100101000000" when "1010101101",
      "1010101110000000000000000001110010111001000011111101101110001001111111100001011" when "1010101110",
      "1010101111000000000000000001110011001110100000111101101110000001001011110000100" when "1010101111",
      "1010110000000000000000000001110011100011111111111101101101111000011001010101100" when "1010110000",
      "1010110001000000000000000001110011111001100000111101101101101111101000010000100" when "1010110001",
      "1010110010000000000000000001110100001111000011111101101101100110111000100001110" when "1010110010",
      "1010110011000000000000000001110100100100101000111101101101011110001010001001001" when "1010110011",
      "1010110100000000000000000001110100111010001111111101101101010101011101000110111" when "1010110100",
      "1010110101000000000000000001110101001111111000111101101101001100110001011011001" when "1010110101",
      "1010110110000000000000000001110101100101100011111101101101000100000111000110000" when "1010110110",
      "1010110111000000000000000001110101111011010000111101101100111011011110000111101" when "1010110111",
      "1010111000000000000000000001110110010000111111111101101100110010110110100000001" when "1010111000",
      "1010111001000000000000000001110110100110110000111101101100101010010000001111110" when "1010111001",
      "1010111010000000000000000001110110111100100011111101101100100001101011010110011" when "1010111010",
      "1010111011000000000000000001110111010010011000111101101100011001000111110100010" when "1010111011",
      "1010111100000000000000000001110111101000001111111101101100010000100101101001100" when "1010111100",
      "1010111101000000000000000001110111111110001000111101101100001000000100110110010" when "1010111101",
      "1010111110000000000000000001111000010100000011111101101011111111100101011010101" when "1010111110",
      "1010111111000000000000000001111000101010000000111101101011110111000111010110111" when "1010111111",
      "1011000000000000000000000001111000111111111111111101101011101110101010101010111" when "1011000000",
      "1011000001000000000000000001111001010110000000111101101011100110001111010110111" when "1011000001",
      "1011000010000000000000000001111001101100000011111101101011011101110101011011000" when "1011000010",
      "1011000011000000000000000001111010000010001000111101101011010101011100110111011" when "1011000011",
      "1011000100000000000000000001111010011000001111111101101011001101000101101100001" when "1011000100",
      "1011000101000000000000000001111010101110011000111101101011000100101111111001011" when "1011000101",
      "1011000110000000000000000001111011000100100011111101101010111100011011011111011" when "1011000110",
      "1011000111000000000000000001111011011010110000111101101010110100001000011110000" when "1011000111",
      "1011001000000000000000000001111011110000111111111101101010101011110110110101100" when "1011001000",
      "1011001001000000000000000001111100000111010000111101101010100011100110100110000" when "1011001001",
      "1011001010000000000000000001111100011101100011111101101010011011010111101111101" when "1011001010",
      "1011001011000000000000000001111100110011111000111101101010010011001010010010100" when "1011001011",
      "1011001100000000000000000001111101001010001111111101101010001010111110001110110" when "1011001100",
      "1011001101000000000000000001111101100000101000111101101010000010110011100100101" when "1011001101",
      "1011001110000000000000000001111101110111000011111101101001111010101010010100000" when "1011001110",
      "1011001111000000000000000001111110001101100000111101101001110010100010011101001" when "1011001111",
      "1011010000000000000000000001111110100011111111111101101001101010011100000000001" when "1011010000",
      "1011010001000000000000000001111110111010100000111101101001100010010110111101001" when "1011010001",
      "1011010010000000000000000001111111010001000011111101101001011010010011010100010" when "1011010010",
      "1011010011000000000000000001111111100111101000111101101001010010010001000101110" when "1011010011",
      "1011010100000000000000000001111111111110001111111101101001001010010000010001100" when "1011010100",
      "1011010101000000000000000010000000010100111000111101101001000010010000110111110" when "1011010101",
      "1011010110000000000000000010000000101011100011111101101000111010010010111000101" when "1011010110",
      "1011010111000000000000000010000001000010010000111101101000110010010110010100010" when "1011010111",
      "1011011000000000000000000010000001011000111111111101101000101010011011001010110" when "1011011000",
      "1011011001000000000000000010000001101111110000111101101000100010100001011100010" when "1011011001",
      "1011011010000000000000000010000010000110100011111101101000011010101001001001000" when "1011011010",
      "1011011011000000000000000010000010011101011000111101101000010010110010010000111" when "1011011011",
      "1011011100000000000000000010000010110100001111111101101000001010111100110100001" when "1011011100",
      "1011011101000000000000000010000011001011001000111101101000000011001000110010111" when "1011011101",
      "1011011110000000000000000010000011100010000011111101100111111011010110001101010" when "1011011110",
      "1011011111000000000000000010000011111001000000111101100111110011100101000011011" when "1011011111",
      "1011100000000000000000000010000100001111111111111101100111101011110101010101011" when "1011100000",
      "1011100001000000000000000010000100100111000000111101100111100100000111000011100" when "1011100001",
      "1011100010000000000000000010000100111110000011111101100111011100011010001101101" when "1011100010",
      "1011100011000000000000000010000101010101001000111101100111010100101110110100000" when "1011100011",
      "1011100100000000000000000010000101101100001111111101100111001101000100110110110" when "1011100100",
      "1011100101000000000000000010000110000011011000111101100111000101011100010110000" when "1011100101",
      "1011100110000000000000000010000110011010100011111101100110111101110101010001111" when "1011100110",
      "1011100111000000000000000010000110110001110000111101100110110110001111101010101" when "1011100111",
      "1011101000000000000000000010000111001000111111111101100110101110101011100000001" when "1011101000",
      "1011101001000000000000000010000111100000010000111101100110100111001000110010101" when "1011101001",
      "1011101010000000000000000010000111110111100011111101100110011111100111100010010" when "1011101010",
      "1011101011000000000000000010001000001110111000111101100110011000000111101111001" when "1011101011",
      "1011101100000000000000000010001000100110001111111101100110010000101001011001011" when "1011101100",
      "1011101101000000000000000010001000111101101000111101100110001001001100100001001" when "1011101101",
      "1011101110000000000000000010001001010101000011111101100110000001110001000110101" when "1011101110",
      "1011101111000000000000000010001001101100100000111101100101111010010111001001110" when "1011101111",
      "1011110000000000000000000010001010000011111111111101100101110010111110101010110" when "1011110000",
      "1011110001000000000000000010001010011011100000111101100101101011100111101001110" when "1011110001",
      "1011110010000000000000000010001010110011000011111101100101100100010010000110111" when "1011110010",
      "1011110011000000000000000010001011001010101000111101100101011100111110000010010" when "1011110011",
      "1011110100000000000000000010001011100010001111111101100101010101101011011100000" when "1011110100",
      "1011110101000000000000000010001011111001111000111101100101001110011010010100011" when "1011110101",
      "1011110110000000000000000010001100010001100011111101100101000111001010101011010" when "1011110110",
      "1011110111000000000000000010001100101001010000111101100100111111111100100000111" when "1011110111",
      "1011111000000000000000000010001101000000111111111101100100111000101111110101011" when "1011111000",
      "1011111001000000000000000010001101011000110000111101100100110001100100101000111" when "1011111001",
      "1011111010000000000000000010001101110000100011111101100100101010011010111011100" when "1011111010",
      "1011111011000000000000000010001110001000011000111101100100100011010010101101100" when "1011111011",
      "1011111100000000000000000010001110100000001111111101100100011100001011111110110" when "1011111100",
      "1011111101000000000000000010001110111000001000111101100100010101000110101111100" when "1011111101",
      "1011111110000000000000000010001111010000000011111101100100001110000010111111111" when "1011111110",
      "1011111111000000000000000010001111101000000000111101100100000111000000110000000" when "1011111111",
      "1100000000000000000000000010001111111111111111111101100100000000000000000000000" when "1100000000",
      "1100000001000000000000000010010000011000000000111101100011111001000000110000000" when "1100000001",
      "1100000010000000000000000010010000110000000011111101100011110010000011000000010" when "1100000010",
      "1100000011000000000000000010010001001000001000111101100011101011000110110000101" when "1100000011",
      "1100000100000000000000000010010001100000001111111101100011100100001100000001011" when "1100000100",
      "1100000101000000000000000010010001111000011000111101100011011101010010110010101" when "1100000101",
      "1100000110000000000000000010010010010000100011111101100011010110011011000100100" when "1100000110",
      "1100000111000000000000000010010010101000110000111101100011001111100100110111001" when "1100000111",
      "1100001000000000000000000010010011000000111111111101100011001000110000001010101" when "1100001000",
      "1100001001000000000000000010010011011001010000111101100011000001111100111111010" when "1100001001",
      "1100001010000000000000000010010011110001100011111101100010111011001011010100111" when "1100001010",
      "1100001011000000000000000010010100001001111000111101100010110100011011001011110" when "1100001011",
      "1100001100000000000000000010010100100010001111111101100010101101101100100100000" when "1100001100",
      "1100001101000000000000000010010100111010101000111101100010100110111111011101110" when "1100001101",
      "1100001110000000000000000010010101010011000011111101100010100000010011111001001" when "1100001110",
      "1100001111000000000000000010010101101011100000111101100010011001101001110110011" when "1100001111",
      "1100010000000000000000000010010110000011111111111101100010010011000001010101011" when "1100010000",
      "1100010001000000000000000010010110011100100000111101100010001100011010010110011" when "1100010001",
      "1100010010000000000000000010010110110101000011111101100010000101110100111001100" when "1100010010",
      "1100010011000000000000000010010111001101101000111101100001111111010000111110111" when "1100010011",
      "1100010100000000000000000010010111100110001111111101100001111000101110100110101" when "1100010100",
      "1100010101000000000000000010010111111110111000111101100001110010001101110000111" when "1100010101",
      "1100010110000000000000000010011000010111100011111101100001101011101110011101111" when "1100010110",
      "1100010111000000000000000010011000110000010000111101100001100101010000101101100" when "1100010111",
      "1100011000000000000000000010011001001000111111111101100001011110110100100000000" when "1100011000",
      "1100011001000000000000000010011001100001110000111101100001011000011001110101100" when "1100011001",
      "1100011010000000000000000010011001111010100011111101100001010010000000101110001" when "1100011010",
      "1100011011000000000000000010011010010011011000111101100001001011101001001010000" when "1100011011",
      "1100011100000000000000000010011010101100001111111101100001000101010011001001010" when "1100011100",
      "1100011101000000000000000010011011000101001000111101100000111110111110101100001" when "1100011101",
      "1100011110000000000000000010011011011110000011111101100000111000101011110010100" when "1100011110",
      "1100011111000000000000000010011011110111000000111101100000110010011010011100101" when "1100011111",
      "1100100000000000000000000010011100001111111111111101100000101100001010101010101" when "1100100000",
      "1100100001000000000000000010011100101001000000111101100000100101111100011100101" when "1100100001",
      "1100100010000000000000000010011101000010000011111101100000011111101111110010110" when "1100100010",
      "1100100011000000000000000010011101011011001000111101100000011001100100101101010" when "1100100011",
      "1100100100000000000000000010011101110100001111111101100000010011011011001100000" when "1100100100",
      "1100100101000000000000000010011110001101011000111101100000001101010011001111010" when "1100100101",
      "1100100110000000000000000010011110100110100011111101100000000111001100110111001" when "1100100110",
      "1100100111000000000000000010011110111111110000111101100000000001001000000011110" when "1100100111",
      "1100101000000000000000000010011111011000111111111101011111111011000100110101010" when "1100101000",
      "1100101001000000000000000010011111110010010000111101011111110101000011001011110" when "1100101001",
      "1100101010000000000000000010100000001011100011111101011111101111000011000111100" when "1100101010",
      "1100101011000000000000000010100000100100111000111101011111101001000100101000011" when "1100101011",
      "1100101100000000000000000010100000111110001111111101011111100011000111101110101" when "1100101100",
      "1100101101000000000000000010100001010111101000111101011111011101001100011010011" when "1100101101",
      "1100101110000000000000000010100001110001000011111101011111010111010010101011110" when "1100101110",
      "1100101111000000000000000010100010001010100000111101011111010001011010100010111" when "1100101111",
      "1100110000000000000000000010100010100011111111111101011111001011100011111111111" when "1100110000",
      "1100110001000000000000000010100010111101100000111101011111000101101111000011000" when "1100110001",
      "1100110010000000000000000010100011010111000011111101011110111111111011101100001" when "1100110010",
      "1100110011000000000000000010100011110000101000111101011110111010001001111011100" when "1100110011",
      "1100110100000000000000000010100100001010001111111101011110110100011001110001010" when "1100110100",
      "1100110101000000000000000010100100100011111000111101011110101110101011001101100" when "1100110101",
      "1100110110000000000000000010100100111101100011111101011110101000111110010000011" when "1100110110",
      "1100110111000000000000000010100101010111010000111101011110100011010010111010001" when "1100110111",
      "1100111000000000000000000010100101110000111111111101011110011101101001001010101" when "1100111000",
      "1100111001000000000000000010100110001010110000111101011110011000000001000010001" when "1100111001",
      "1100111010000000000000000010100110100100100011111101011110010010011010100000110" when "1100111010",
      "1100111011000000000000000010100110111110011000111101011110001100110101100110101" when "1100111011",
      "1100111100000000000000000010100111011000001111111101011110000111010010010011111" when "1100111100",
      "1100111101000000000000000010100111110010001000111101011110000001110000101000101" when "1100111101",
      "1100111110000000000000000010101000001100000011111101011101111100010000100101001" when "1100111110",
      "1100111111000000000000000010101000100110000000111101011101110110110010001001010" when "1100111111",
      "1101000000000000000000000010101000111111111111111101011101110001010101010101010" when "1101000000",
      "1101000001000000000000000010101001011010000000111101011101101011111010001001010" when "1101000001",
      "1101000010000000000000000010101001110100000011111101011101100110100000100101011" when "1101000010",
      "1101000011000000000000000010101010001110001000111101011101100001001000101001110" when "1101000011",
      "1101000100000000000000000010101010101000001111111101011101011011110010010110100" when "1101000100",
      "1101000101000000000000000010101011000010011000111101011101010110011101101011111" when "1101000101",
      "1101000110000000000000000010101011011100100011111101011101010001001010101001110" when "1101000110",
      "1101000111000000000000000010101011110110110000111101011101001011111001010000011" when "1101000111",
      "1101001000000000000000000010101100010000111111111101011101000110101001011111111" when "1101001000",
      "1101001001000000000000000010101100101011010000111101011101000001011011011000011" when "1101001001",
      "1101001010000000000000000010101101000101100011111101011100111100001110111010000" when "1101001010",
      "1101001011000000000000000010101101011111111000111101011100110111000100000100111" when "1101001011",
      "1101001100000000000000000010101101111010001111111101011100110001111010111001010" when "1101001100",
      "1101001101000000000000000010101110010100101000111101011100101100110011010111000" when "1101001101",
      "1101001110000000000000000010101110101111000011111101011100100111101101011110011" when "1101001110",
      "1101001111000000000000000010101111001001100000111101011100100010101001001111100" when "1101001111",
      "1101010000000000000000000010101111100011111111111101011100011101100110101010100" when "1101010000",
      "1101010001000000000000000010101111111110100000111101011100011000100101101111100" when "1101010001",
      "1101010010000000000000000010110000011001000011111101011100010011100110011110110" when "1101010010",
      "1101010011000000000000000010110000110011101000111101011100001110101000111000001" when "1101010011",
      "1101010100000000000000000010110001001110001111111101011100001001101100111011111" when "1101010100",
      "1101010101000000000000000010110001101000111000111101011100000100110010101010001" when "1101010101",
      "1101010110000000000000000010110010000011100011111101011011111111111010000011000" when "1101010110",
      "1101010111000000000000000010110010011110010000111101011011111011000011000110101" when "1101010111",
      "1101011000000000000000000010110010111000111111111101011011110110001101110101001" when "1101011000",
      "1101011001000000000000000010110011010011110000111101011011110001011010001110110" when "1101011001",
      "1101011010000000000000000010110011101110100011111101011011101100101000010011011" when "1101011010",
      "1101011011000000000000000010110100001001011000111101011011100111111000000011010" when "1101011011",
      "1101011100000000000000000010110100100100001111111101011011100011001001011110100" when "1101011100",
      "1101011101000000000000000010110100111111001000111101011011011110011100100101010" when "1101011101",
      "1101011110000000000000000010110101011010000011111101011011011001110001010111101" when "1101011110",
      "1101011111000000000000000010110101110101000000111101011011010101000111110101110" when "1101011111",
      "1101100000000000000000000010110110001111111111111101011011010000011111111111111" when "1101100000",
      "1101100001000000000000000010110110101011000000111101011011001011111001110101111" when "1101100001",
      "1101100010000000000000000010110111000110000011111101011011000111010101011000000" when "1101100010",
      "1101100011000000000000000010110111100001001000111101011011000010110010100110011" when "1101100011",
      "1101100100000000000000000010110111111100001111111101011010111110010001100001001" when "1101100100",
      "1101100101000000000000000010111000010111011000111101011010111001110010001000011" when "1101100101",
      "1101100110000000000000000010111000110010100011111101011010110101010100011100011" when "1101100110",
      "1101100111000000000000000010111001001101110000111101011010110000111000011101000" when "1101100111",
      "1101101000000000000000000010111001101000111111111101011010101100011110001010100" when "1101101000",
      "1101101001000000000000000010111010000100010000111101011010101000000101100101000" when "1101101001",
      "1101101010000000000000000010111010011111100011111101011010100011101110101100101" when "1101101010",
      "1101101011000000000000000010111010111010111000111101011010011111011001100001100" when "1101101011",
      "1101101100000000000000000010111011010110001111111101011010011011000110000011110" when "1101101100",
      "1101101101000000000000000010111011110001101000111101011010010110110100010011101" when "1101101101",
      "1101101110000000000000000010111100001101000011111101011010010010100100010001000" when "1101101110",
      "1101101111000000000000000010111100101000100000111101011010001110010101111100001" when "1101101111",
      "1101110000000000000000000010111101000011111111111101011010001010001001010101001" when "1101110000",
      "1101110001000000000000000010111101011111100000111101011010000101111110011100001" when "1101110001",
      "1101110010000000000000000010111101111011000011111101011010000001110101010001010" when "1101110010",
      "1101110011000000000000000010111110010110101000111101011001111101101101110100101" when "1101110011",
      "1101110100000000000000000010111110110010001111111101011001111001101000000110100" when "1101110100",
      "1101110101000000000000000010111111001101111000111101011001110101100100000110110" when "1101110101",
      "1101110110000000000000000010111111101001100011111101011001110001100001110101101" when "1101110110",
      "1101110111000000000000000011000000000101010000111101011001101101100001010011010" when "1101110111",
      "1101111000000000000000000011000000100000111111111101011001101001100010011111110" when "1101111000",
      "1101111001000000000000000011000000111100110000111101011001100101100101011011010" when "1101111001",
      "1101111010000000000000000011000001011000100011111101011001100001101010000110000" when "1101111010",
      "1101111011000000000000000011000001110100011000111101011001011101110000011111111" when "1101111011",
      "1101111100000000000000000011000010010000001111111101011001011001111000101001001" when "1101111100",
      "1101111101000000000000000011000010101100001000111101011001010110000010100001111" when "1101111101",
      "1101111110000000000000000011000011001000000011111101011001010010001110001010010" when "1101111110",
      "1101111111000000000000000011000011100100000000111101011001001110011011100010011" when "1101111111",
      "1110000000000000000000000011000011111111111111111101011001001010101010101010011" when "1110000000",
      "1110000001000000000000000011000100011100000000111101011001000110111011100010100" when "1110000001",
      "1110000010000000000000000011000100111000000011111101011001000011001110001010101" when "1110000010",
      "1110000011000000000000000011000101010100001000111101011000111111100010100011000" when "1110000011",
      "1110000100000000000000000011000101110000001111111101011000111011111000101011110" when "1110000100",
      "1110000101000000000000000011000110001100011000111101011000111000010000100101000" when "1110000101",
      "1110000110000000000000000011000110101000100011111101011000110100101010001110111" when "1110000110",
      "1110000111000000000000000011000111000100110000111101011000110001000101101001100" when "1110000111",
      "1110001000000000000000000011000111100000111111111101011000101101100010110101001" when "1110001000",
      "1110001001000000000000000011000111111101010000111101011000101010000001110001101" when "1110001001",
      "1110001010000000000000000011001000011001100011111101011000100110100010011111010" when "1110001010",
      "1110001011000000000000000011001000110101111000111101011000100011000100111110001" when "1110001011",
      "1110001100000000000000000011001001010010001111111101011000011111101001001110011" when "1110001100",
      "1110001101000000000000000011001001101110101000111101011000011100001111010000001" when "1110001101",
      "1110001110000000000000000011001010001011000011111101011000011000110111000011101" when "1110001110",
      "1110001111000000000000000011001010100111100000111101011000010101100000101000110" when "1110001111",
      "1110010000000000000000000011001011000011111111111101011000010010001011111111110" when "1110010000",
      "1110010001000000000000000011001011100000100000111101011000001110111001001000110" when "1110010001",
      "1110010010000000000000000011001011111101000011111101011000001011101000000011111" when "1110010010",
      "1110010011000000000000000011001100011001101000111101011000001000011000110001010" when "1110010011",
      "1110010100000000000000000011001100110110001111111101011000000101001011010001000" when "1110010100",
      "1110010101000000000000000011001101010010111000111101011000000001111111100011011" when "1110010101",
      "1110010110000000000000000011001101101111100011111101010111111110110101101000010" when "1110010110",
      "1110010111000000000000000011001110001100010000111101010111111011101101011111111" when "1110010111",
      "1110011000000000000000000011001110101000111111111101010111111000100111001010011" when "1110011000",
      "1110011001000000000000000011001111000101110000111101010111110101100010100111111" when "1110011001",
      "1110011010000000000000000011001111100010100011111101010111110010011111111000100" when "1110011010",
      "1110011011000000000000000011001111111111011000111101010111101111011110111100011" when "1110011011",
      "1110011100000000000000000011010000011100001111111101010111101100011111110011110" when "1110011100",
      "1110011101000000000000000011010000111001001000111101010111101001100010011110100" when "1110011101",
      "1110011110000000000000000011010001010110000011111101010111100110100110111100111" when "1110011110",
      "1110011111000000000000000011010001110011000000111101010111100011101101001111000" when "1110011111",
      "1110100000000000000000000011010010001111111111111101010111100000110101010101000" when "1110100000",
      "1110100001000000000000000011010010101101000000111101010111011101111111001111000" when "1110100001",
      "1110100010000000000000000011010011001010000011111101010111011011001010111101010" when "1110100010",
      "1110100011000000000000000011010011100111001000111101010111011000011000011111101" when "1110100011",
      "1110100100000000000000000011010100000100001111111101010111010101100111110110011" when "1110100100",
      "1110100101000000000000000011010100100001011000111101010111010010111001000001101" when "1110100101",
      "1110100110000000000000000011010100111110100011111101010111010000001100000001100" when "1110100110",
      "1110100111000000000000000011010101011011110000111101010111001101100000110110001" when "1110100111",
      "1110101000000000000000000011010101111000111111111101010111001010110111011111101" when "1110101000",
      "1110101001000000000000000011010110010110010000111101010111001000001111111110010" when "1110101001",
      "1110101010000000000000000011010110110011100011111101010111000101101010010001111" when "1110101010",
      "1110101011000000000000000011010111010000111000111101010111000011000110011010110" when "1110101011",
      "1110101100000000000000000011010111101110001111111101010111000000100100011001000" when "1110101100",
      "1110101101000000000000000011011000001011101000111101010110111110000100001100110" when "1110101101",
      "1110101110000000000000000011011000101001000011111101010110111011100101110110001" when "1110101110",
      "1110101111000000000000000011011001000110100000111101010110111001001001010101010" when "1110101111",
      "1110110000000000000000000011011001100011111111111101010110110110101110101010011" when "1110110000",
      "1110110001000000000000000011011010000001100000111101010110110100010101110101011" when "1110110001",
      "1110110010000000000000000011011010011111000011111101010110110001111110110110100" when "1110110010",
      "1110110011000000000000000011011010111100101000111101010110101111101001101101111" when "1110110011",
      "1110110100000000000000000011011011011010001111111101010110101101010110011011101" when "1110110100",
      "1110110101000000000000000011011011110111111000111101010110101011000100111111111" when "1110110101",
      "1110110110000000000000000011011100010101100011111101010110101000110101011010111" when "1110110110",
      "1110110111000000000000000011011100110011010000111101010110100110100111101100100" when "1110110111",
      "1110111000000000000000000011011101010000111111111101010110100100011011110101000" when "1110111000",
      "1110111001000000000000000011011101101110110000111101010110100010010001110100100" when "1110111001",
      "1110111010000000000000000011011110001100100011111101010110100000001001101011001" when "1110111010",
      "1110111011000000000000000011011110101010011000111101010110011110000011011001000" when "1110111011",
      "1110111100000000000000000011011111001000001111111101010110011011111110111110010" when "1110111100",
      "1110111101000000000000000011011111100110001000111101010110011001111100011011001" when "1110111101",
      "1110111110000000000000000011100000000100000011111101010110010111111011101111100" when "1110111110",
      "1110111111000000000000000011100000100010000000111101010110010101111100111011101" when "1110111111",
      "1111000000000000000000000011100000111111111111111101010110010011111111111111101" when "1111000000",
      "1111000001000000000000000011100001011110000000111101010110010010000100111011101" when "1111000001",
      "1111000010000000000000000011100001111100000011111101010110010000001011101111110" when "1111000010",
      "1111000011000000000000000011100010011010001000111101010110001110010100011100001" when "1111000011",
      "1111000100000000000000000011100010111000001111111101010110001100011111000001000" when "1111000100",
      "1111000101000000000000000011100011010110011000111101010110001010101011011110010" when "1111000101",
      "1111000110000000000000000011100011110100100011111101010110001000111001110100001" when "1111000110",
      "1111000111000000000000000011100100010010110000111101010110000111001010000010110" when "1111000111",
      "1111001000000000000000000011100100110000111111111101010110000101011100001010010" when "1111001000",
      "1111001001000000000000000011100101001111010000111101010110000011110000001010110" when "1111001001",
      "1111001010000000000000000011100101101101100011111101010110000010000110000100100" when "1111001010",
      "1111001011000000000000000011100110001011111000111101010110000000011101110111011" when "1111001011",
      "1111001100000000000000000011100110101010001111111101010101111110110111100011101" when "1111001100",
      "1111001101000000000000000011100111001000101000111101010101111101010011001001011" when "1111001101",
      "1111001110000000000000000011100111100111000011111101010101111011110000101000110" when "1111001110",
      "1111001111000000000000000011101000000101100000111101010101111010010000000001111" when "1111001111",
      "1111010000000000000000000011101000100011111111111101010101111000110001010100111" when "1111010000",
      "1111010001000000000000000011101001000010100000111101010101110111010100100010000" when "1111010001",
      "1111010010000000000000000011101001100001000011111101010101110101111001101001001" when "1111010010",
      "1111010011000000000000000011101001111111101000111101010101110100100000101010100" when "1111010011",
      "1111010100000000000000000011101010011110001111111101010101110011001001100110010" when "1111010100",
      "1111010101000000000000000011101010111100111000111101010101110001110100011100100" when "1111010101",
      "1111010110000000000000000011101011011011100011111101010101110000100001001101011" when "1111010110",
      "1111010111000000000000000011101011111010010000111101010101101111001111111001000" when "1111010111",
      "1111011000000000000000000011101100011000111111111101010101101110000000011111101" when "1111011000",
      "1111011001000000000000000011101100110111110000111101010101101100110011000001001" when "1111011001",
      "1111011010000000000000000011101101010110100011111101010101101011100111011101110" when "1111011010",
      "1111011011000000000000000011101101110101011000111101010101101010011101110101101" when "1111011011",
      "1111011100000000000000000011101110010100001111111101010101101001010110001000111" when "1111011100",
      "1111011101000000000000000011101110110011001000111101010101101000010000010111101" when "1111011101",
      "1111011110000000000000000011101111010010000011111101010101100111001100100010001" when "1111011110",
      "1111011111000000000000000011101111110001000000111101010101100110001010101000010" when "1111011111",
      "1111100000000000000000000011110000001111111111111101010101100101001010101010010" when "1111100000",
      "1111100001000000000000000011110000101111000000111101010101100100001100101000010" when "1111100001",
      "1111100010000000000000000011110001001110000011111101010101100011010000100010011" when "1111100010",
      "1111100011000000000000000011110001101101001000111101010101100010010110011000110" when "1111100011",
      "1111100100000000000000000011110010001100001111111101010101100001011110001011100" when "1111100100",
      "1111100101000000000000000011110010101011011000111101010101100000100111111010111" when "1111100101",
      "1111100110000000000000000011110011001010100011111101010101011111110011100110110" when "1111100110",
      "1111100111000000000000000011110011101001110000111101010101011111000001001111011" when "1111100111",
      "1111101000000000000000000011110100001000111111111101010101011110010000110100111" when "1111101000",
      "1111101001000000000000000011110100101000010000111101010101011101100010010111011" when "1111101001",
      "1111101010000000000000000011110101000111100011111101010101011100110101110111000" when "1111101010",
      "1111101011000000000000000011110101100110111000111101010101011100001011010011111" when "1111101011",
      "1111101100000000000000000011110110000110001111111101010101011011100010101110010" when "1111101100",
      "1111101101000000000000000011110110100101101000111101010101011010111100000110000" when "1111101101",
      "1111101110000000000000000011110111000101000011111101010101011010010111011011011" when "1111101110",
      "1111101111000000000000000011110111100100100000111101010101011001110100101110100" when "1111101111",
      "1111110000000000000000000011111000000011111111111101010101011001010011111111100" when "1111110000",
      "1111110001000000000000000011111000100011100000111101010101011000110101001110100" when "1111110001",
      "1111110010000000000000000011111001000011000011111101010101011000011000011011110" when "1111110010",
      "1111110011000000000000000011111001100010101000111101010101010111111101100111001" when "1111110011",
      "1111110100000000000000000011111010000010001111111101010101010111100100110000111" when "1111110100",
      "1111110101000000000000000011111010100001111000111101010101010111001101111001001" when "1111110101",
      "1111110110000000000000000011111011000001100011111101010101010110111001000000000" when "1111110110",
      "1111110111000000000000000011111011100001010000111101010101010110100110000101101" when "1111110111",
      "1111111000000000000000000011111100000000111111111101010101010110010101001010001" when "1111111000",
      "1111111001000000000000000011111100100000110000111101010101010110000110001101110" when "1111111001",
      "1111111010000000000000000011111101000000100011111101010101010101111001010000011" when "1111111010",
      "1111111011000000000000000011111101100000011000111101010101010101101110010010010" when "1111111011",
      "1111111100000000000000000011111110000000001111111101010101010101100101010011100" when "1111111100",
      "1111111101000000000000000011111110100000001000111101010101010101011110010100010" when "1111111101",
      "1111111110000000000000000011111111000000000011111101010101010101011001010100101" when "1111111110",
      "1111111111000000000000000011111111100000000000111101010101010101010110010100111" when "1111111111",
      "-------------------------------------------------------------------------------" when others;
   Y1_c5 <= Y0_c5; -- for the possible blockram register
   Y <= Y1_c5;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_104_Freq300_uid53
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_104_Freq300_uid53 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(103 downto 0);
          Y : in  std_logic_vector(103 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(103 downto 0)   );
end entity;

architecture arch of IntAdder_104_Freq300_uid53 is
signal Rtmp_c6 :  std_logic_vector(103 downto 0);
signal X_c5, X_c6 :  std_logic_vector(103 downto 0);
signal Y_c6 :  std_logic_vector(103 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               X_c5 <= X;
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
               Y_c6 <= Y;
               Cin_c6 <= Cin_c5;
            end if;
         end if;
      end process;
   Rtmp_c6 <= X_c6 + Y_c6 + Cin_c6;
   R <= Rtmp_c6;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_104_Freq300_uid56
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_104_Freq300_uid56 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(103 downto 0);
          Y : in  std_logic_vector(103 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(103 downto 0)   );
end entity;

architecture arch of IntAdder_104_Freq300_uid56 is
signal Rtmp_c8 :  std_logic_vector(103 downto 0);
signal X_c7, X_c8 :  std_logic_vector(103 downto 0);
signal Y_c8 :  std_logic_vector(103 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               X_c7 <= X;
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
               Y_c8 <= Y;
               Cin_c8 <= Cin_c7;
            end if;
         end if;
      end process;
   Rtmp_c8 <= X_c8 + Y_c8 + Cin_c8;
   R <= Rtmp_c8;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_82_Freq300_uid68
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_82_Freq300_uid68 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(81 downto 0);
          Y : in  std_logic_vector(81 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(81 downto 0)   );
end entity;

architecture arch of IntAdder_82_Freq300_uid68 is
signal Cin_1_c0, Cin_1_c1 :  std_logic;
signal X_1_c0, X_1_c1 :  std_logic_vector(82 downto 0);
signal Y_1_c0, Y_1_c1 :  std_logic_vector(82 downto 0);
signal S_1_c1 :  std_logic_vector(82 downto 0);
signal R_1_c1 :  std_logic_vector(81 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_1_c1 <= Cin_1_c0;
               X_1_c1 <= X_1_c0;
               Y_1_c1 <= Y_1_c0;
            end if;
         end if;
      end process;
   Cin_1_c0 <= Cin;
   X_1_c0 <= '0' & X(81 downto 0);
   Y_1_c0 <= '0' & Y(81 downto 0);
   S_1_c1 <= X_1_c1 + Y_1_c1 + Cin_1_c1;
   R_1_c1 <= S_1_c1(81 downto 0);
   R <= R_1_c1 ;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq300_uid58
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid58 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          R : out  std_logic_vector(80 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid58 is
   component FixRealKCM_Freq300_uid58_T0_Freq300_uid61 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(80 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid58_T1_Freq300_uid64 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(75 downto 0)   );
   end component;

   component IntAdder_82_Freq300_uid68 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(81 downto 0);
             Y : in  std_logic_vector(81 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(81 downto 0)   );
   end component;

signal FixRealKCM_Freq300_uid58_A0_c0 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid58_T0_c0 :  std_logic_vector(80 downto 0);
signal FixRealKCM_Freq300_uid58_T0_copy62_c0 :  std_logic_vector(80 downto 0);
signal bh59_w0_0_c0 :  std_logic;
signal bh59_w1_0_c0 :  std_logic;
signal bh59_w2_0_c0 :  std_logic;
signal bh59_w3_0_c0 :  std_logic;
signal bh59_w4_0_c0 :  std_logic;
signal bh59_w5_0_c0 :  std_logic;
signal bh59_w6_0_c0 :  std_logic;
signal bh59_w7_0_c0 :  std_logic;
signal bh59_w8_0_c0 :  std_logic;
signal bh59_w9_0_c0 :  std_logic;
signal bh59_w10_0_c0 :  std_logic;
signal bh59_w11_0_c0 :  std_logic;
signal bh59_w12_0_c0 :  std_logic;
signal bh59_w13_0_c0 :  std_logic;
signal bh59_w14_0_c0 :  std_logic;
signal bh59_w15_0_c0 :  std_logic;
signal bh59_w16_0_c0 :  std_logic;
signal bh59_w17_0_c0 :  std_logic;
signal bh59_w18_0_c0 :  std_logic;
signal bh59_w19_0_c0 :  std_logic;
signal bh59_w20_0_c0 :  std_logic;
signal bh59_w21_0_c0 :  std_logic;
signal bh59_w22_0_c0 :  std_logic;
signal bh59_w23_0_c0 :  std_logic;
signal bh59_w24_0_c0 :  std_logic;
signal bh59_w25_0_c0 :  std_logic;
signal bh59_w26_0_c0 :  std_logic;
signal bh59_w27_0_c0 :  std_logic;
signal bh59_w28_0_c0 :  std_logic;
signal bh59_w29_0_c0 :  std_logic;
signal bh59_w30_0_c0 :  std_logic;
signal bh59_w31_0_c0 :  std_logic;
signal bh59_w32_0_c0 :  std_logic;
signal bh59_w33_0_c0 :  std_logic;
signal bh59_w34_0_c0 :  std_logic;
signal bh59_w35_0_c0 :  std_logic;
signal bh59_w36_0_c0 :  std_logic;
signal bh59_w37_0_c0 :  std_logic;
signal bh59_w38_0_c0 :  std_logic;
signal bh59_w39_0_c0 :  std_logic;
signal bh59_w40_0_c0 :  std_logic;
signal bh59_w41_0_c0 :  std_logic;
signal bh59_w42_0_c0 :  std_logic;
signal bh59_w43_0_c0 :  std_logic;
signal bh59_w44_0_c0 :  std_logic;
signal bh59_w45_0_c0 :  std_logic;
signal bh59_w46_0_c0 :  std_logic;
signal bh59_w47_0_c0 :  std_logic;
signal bh59_w48_0_c0 :  std_logic;
signal bh59_w49_0_c0 :  std_logic;
signal bh59_w50_0_c0 :  std_logic;
signal bh59_w51_0_c0 :  std_logic;
signal bh59_w52_0_c0 :  std_logic;
signal bh59_w53_0_c0 :  std_logic;
signal bh59_w54_0_c0 :  std_logic;
signal bh59_w55_0_c0 :  std_logic;
signal bh59_w56_0_c0 :  std_logic;
signal bh59_w57_0_c0 :  std_logic;
signal bh59_w58_0_c0 :  std_logic;
signal bh59_w59_0_c0 :  std_logic;
signal bh59_w60_0_c0 :  std_logic;
signal bh59_w61_0_c0 :  std_logic;
signal bh59_w62_0_c0 :  std_logic;
signal bh59_w63_0_c0 :  std_logic;
signal bh59_w64_0_c0 :  std_logic;
signal bh59_w65_0_c0 :  std_logic;
signal bh59_w66_0_c0 :  std_logic;
signal bh59_w67_0_c0 :  std_logic;
signal bh59_w68_0_c0 :  std_logic;
signal bh59_w69_0_c0 :  std_logic;
signal bh59_w70_0_c0 :  std_logic;
signal bh59_w71_0_c0 :  std_logic;
signal bh59_w72_0_c0 :  std_logic;
signal bh59_w73_0_c0 :  std_logic;
signal bh59_w74_0_c0 :  std_logic;
signal bh59_w75_0_c0 :  std_logic;
signal bh59_w76_0_c0 :  std_logic;
signal bh59_w77_0_c0 :  std_logic;
signal bh59_w78_0_c0 :  std_logic;
signal bh59_w79_0_c0 :  std_logic;
signal bh59_w80_0_c0 :  std_logic;
signal FixRealKCM_Freq300_uid58_A1_c0 :  std_logic_vector(5 downto 0);
signal FixRealKCM_Freq300_uid58_T1_c0 :  std_logic_vector(75 downto 0);
signal FixRealKCM_Freq300_uid58_T1_copy65_c0 :  std_logic_vector(75 downto 0);
signal bh59_w0_1_c0 :  std_logic;
signal bh59_w1_1_c0 :  std_logic;
signal bh59_w2_1_c0 :  std_logic;
signal bh59_w3_1_c0 :  std_logic;
signal bh59_w4_1_c0 :  std_logic;
signal bh59_w5_1_c0 :  std_logic;
signal bh59_w6_1_c0 :  std_logic;
signal bh59_w7_1_c0 :  std_logic;
signal bh59_w8_1_c0 :  std_logic;
signal bh59_w9_1_c0 :  std_logic;
signal bh59_w10_1_c0 :  std_logic;
signal bh59_w11_1_c0 :  std_logic;
signal bh59_w12_1_c0 :  std_logic;
signal bh59_w13_1_c0 :  std_logic;
signal bh59_w14_1_c0 :  std_logic;
signal bh59_w15_1_c0 :  std_logic;
signal bh59_w16_1_c0 :  std_logic;
signal bh59_w17_1_c0 :  std_logic;
signal bh59_w18_1_c0 :  std_logic;
signal bh59_w19_1_c0 :  std_logic;
signal bh59_w20_1_c0 :  std_logic;
signal bh59_w21_1_c0 :  std_logic;
signal bh59_w22_1_c0 :  std_logic;
signal bh59_w23_1_c0 :  std_logic;
signal bh59_w24_1_c0 :  std_logic;
signal bh59_w25_1_c0 :  std_logic;
signal bh59_w26_1_c0 :  std_logic;
signal bh59_w27_1_c0 :  std_logic;
signal bh59_w28_1_c0 :  std_logic;
signal bh59_w29_1_c0 :  std_logic;
signal bh59_w30_1_c0 :  std_logic;
signal bh59_w31_1_c0 :  std_logic;
signal bh59_w32_1_c0 :  std_logic;
signal bh59_w33_1_c0 :  std_logic;
signal bh59_w34_1_c0 :  std_logic;
signal bh59_w35_1_c0 :  std_logic;
signal bh59_w36_1_c0 :  std_logic;
signal bh59_w37_1_c0 :  std_logic;
signal bh59_w38_1_c0 :  std_logic;
signal bh59_w39_1_c0 :  std_logic;
signal bh59_w40_1_c0 :  std_logic;
signal bh59_w41_1_c0 :  std_logic;
signal bh59_w42_1_c0 :  std_logic;
signal bh59_w43_1_c0 :  std_logic;
signal bh59_w44_1_c0 :  std_logic;
signal bh59_w45_1_c0 :  std_logic;
signal bh59_w46_1_c0 :  std_logic;
signal bh59_w47_1_c0 :  std_logic;
signal bh59_w48_1_c0 :  std_logic;
signal bh59_w49_1_c0 :  std_logic;
signal bh59_w50_1_c0 :  std_logic;
signal bh59_w51_1_c0 :  std_logic;
signal bh59_w52_1_c0 :  std_logic;
signal bh59_w53_1_c0 :  std_logic;
signal bh59_w54_1_c0 :  std_logic;
signal bh59_w55_1_c0 :  std_logic;
signal bh59_w56_1_c0 :  std_logic;
signal bh59_w57_1_c0 :  std_logic;
signal bh59_w58_1_c0 :  std_logic;
signal bh59_w59_1_c0 :  std_logic;
signal bh59_w60_1_c0 :  std_logic;
signal bh59_w61_1_c0 :  std_logic;
signal bh59_w62_1_c0 :  std_logic;
signal bh59_w63_1_c0 :  std_logic;
signal bh59_w64_1_c0 :  std_logic;
signal bh59_w65_1_c0 :  std_logic;
signal bh59_w66_1_c0 :  std_logic;
signal bh59_w67_1_c0 :  std_logic;
signal bh59_w68_1_c0 :  std_logic;
signal bh59_w69_1_c0 :  std_logic;
signal bh59_w70_1_c0 :  std_logic;
signal bh59_w71_1_c0 :  std_logic;
signal bh59_w72_1_c0 :  std_logic;
signal bh59_w73_1_c0 :  std_logic;
signal bh59_w74_1_c0 :  std_logic;
signal bh59_w75_1_c0 :  std_logic;
signal bitheapFinalAdd_bh59_In0_c0 :  std_logic_vector(81 downto 0);
signal bitheapFinalAdd_bh59_In1_c0 :  std_logic_vector(81 downto 0);
signal bitheapFinalAdd_bh59_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh59_Out_c1 :  std_logic_vector(81 downto 0);
signal bitheapResult_bh59_c1 :  std_logic_vector(80 downto 0);
signal OutRes_c1 :  std_logic_vector(80 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
            end if;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq300_uid58_A0_c0 <= X(10 downto 6);-- input address  m=10  l=6
   FixRealKCM_Freq300_uid58_Table0: FixRealKCM_Freq300_uid58_T0_Freq300_uid61
      port map ( X => FixRealKCM_Freq300_uid58_A0_c0,
                 Y => FixRealKCM_Freq300_uid58_T0_copy62_c0);
   FixRealKCM_Freq300_uid58_T0_c0 <= FixRealKCM_Freq300_uid58_T0_copy62_c0; -- output copy to hold a pipeline register if needed
   bh59_w0_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(0);
   bh59_w1_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(1);
   bh59_w2_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(2);
   bh59_w3_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(3);
   bh59_w4_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(4);
   bh59_w5_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(5);
   bh59_w6_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(6);
   bh59_w7_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(7);
   bh59_w8_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(8);
   bh59_w9_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(9);
   bh59_w10_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(10);
   bh59_w11_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(11);
   bh59_w12_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(12);
   bh59_w13_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(13);
   bh59_w14_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(14);
   bh59_w15_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(15);
   bh59_w16_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(16);
   bh59_w17_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(17);
   bh59_w18_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(18);
   bh59_w19_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(19);
   bh59_w20_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(20);
   bh59_w21_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(21);
   bh59_w22_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(22);
   bh59_w23_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(23);
   bh59_w24_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(24);
   bh59_w25_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(25);
   bh59_w26_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(26);
   bh59_w27_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(27);
   bh59_w28_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(28);
   bh59_w29_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(29);
   bh59_w30_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(30);
   bh59_w31_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(31);
   bh59_w32_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(32);
   bh59_w33_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(33);
   bh59_w34_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(34);
   bh59_w35_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(35);
   bh59_w36_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(36);
   bh59_w37_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(37);
   bh59_w38_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(38);
   bh59_w39_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(39);
   bh59_w40_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(40);
   bh59_w41_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(41);
   bh59_w42_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(42);
   bh59_w43_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(43);
   bh59_w44_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(44);
   bh59_w45_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(45);
   bh59_w46_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(46);
   bh59_w47_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(47);
   bh59_w48_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(48);
   bh59_w49_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(49);
   bh59_w50_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(50);
   bh59_w51_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(51);
   bh59_w52_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(52);
   bh59_w53_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(53);
   bh59_w54_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(54);
   bh59_w55_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(55);
   bh59_w56_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(56);
   bh59_w57_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(57);
   bh59_w58_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(58);
   bh59_w59_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(59);
   bh59_w60_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(60);
   bh59_w61_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(61);
   bh59_w62_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(62);
   bh59_w63_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(63);
   bh59_w64_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(64);
   bh59_w65_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(65);
   bh59_w66_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(66);
   bh59_w67_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(67);
   bh59_w68_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(68);
   bh59_w69_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(69);
   bh59_w70_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(70);
   bh59_w71_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(71);
   bh59_w72_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(72);
   bh59_w73_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(73);
   bh59_w74_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(74);
   bh59_w75_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(75);
   bh59_w76_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(76);
   bh59_w77_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(77);
   bh59_w78_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(78);
   bh59_w79_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(79);
   bh59_w80_0_c0 <= FixRealKCM_Freq300_uid58_T0_c0(80);
   FixRealKCM_Freq300_uid58_A1_c0 <= X(5 downto 0);-- input address  m=5  l=0
   FixRealKCM_Freq300_uid58_Table1: FixRealKCM_Freq300_uid58_T1_Freq300_uid64
      port map ( X => FixRealKCM_Freq300_uid58_A1_c0,
                 Y => FixRealKCM_Freq300_uid58_T1_copy65_c0);
   FixRealKCM_Freq300_uid58_T1_c0 <= FixRealKCM_Freq300_uid58_T1_copy65_c0; -- output copy to hold a pipeline register if needed
   bh59_w0_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(0);
   bh59_w1_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(1);
   bh59_w2_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(2);
   bh59_w3_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(3);
   bh59_w4_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(4);
   bh59_w5_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(5);
   bh59_w6_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(6);
   bh59_w7_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(7);
   bh59_w8_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(8);
   bh59_w9_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(9);
   bh59_w10_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(10);
   bh59_w11_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(11);
   bh59_w12_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(12);
   bh59_w13_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(13);
   bh59_w14_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(14);
   bh59_w15_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(15);
   bh59_w16_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(16);
   bh59_w17_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(17);
   bh59_w18_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(18);
   bh59_w19_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(19);
   bh59_w20_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(20);
   bh59_w21_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(21);
   bh59_w22_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(22);
   bh59_w23_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(23);
   bh59_w24_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(24);
   bh59_w25_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(25);
   bh59_w26_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(26);
   bh59_w27_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(27);
   bh59_w28_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(28);
   bh59_w29_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(29);
   bh59_w30_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(30);
   bh59_w31_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(31);
   bh59_w32_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(32);
   bh59_w33_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(33);
   bh59_w34_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(34);
   bh59_w35_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(35);
   bh59_w36_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(36);
   bh59_w37_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(37);
   bh59_w38_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(38);
   bh59_w39_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(39);
   bh59_w40_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(40);
   bh59_w41_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(41);
   bh59_w42_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(42);
   bh59_w43_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(43);
   bh59_w44_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(44);
   bh59_w45_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(45);
   bh59_w46_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(46);
   bh59_w47_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(47);
   bh59_w48_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(48);
   bh59_w49_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(49);
   bh59_w50_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(50);
   bh59_w51_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(51);
   bh59_w52_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(52);
   bh59_w53_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(53);
   bh59_w54_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(54);
   bh59_w55_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(55);
   bh59_w56_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(56);
   bh59_w57_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(57);
   bh59_w58_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(58);
   bh59_w59_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(59);
   bh59_w60_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(60);
   bh59_w61_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(61);
   bh59_w62_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(62);
   bh59_w63_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(63);
   bh59_w64_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(64);
   bh59_w65_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(65);
   bh59_w66_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(66);
   bh59_w67_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(67);
   bh59_w68_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(68);
   bh59_w69_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(69);
   bh59_w70_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(70);
   bh59_w71_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(71);
   bh59_w72_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(72);
   bh59_w73_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(73);
   bh59_w74_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(74);
   bh59_w75_1_c0 <= FixRealKCM_Freq300_uid58_T1_c0(75);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh59_In0_c0 <= "0" & bh59_w80_0_c0 & bh59_w79_0_c0 & bh59_w78_0_c0 & bh59_w77_0_c0 & bh59_w76_0_c0 & bh59_w75_0_c0 & bh59_w74_0_c0 & bh59_w73_0_c0 & bh59_w72_0_c0 & bh59_w71_0_c0 & bh59_w70_0_c0 & bh59_w69_0_c0 & bh59_w68_0_c0 & bh59_w67_0_c0 & bh59_w66_0_c0 & bh59_w65_0_c0 & bh59_w64_0_c0 & bh59_w63_0_c0 & bh59_w62_0_c0 & bh59_w61_0_c0 & bh59_w60_0_c0 & bh59_w59_0_c0 & bh59_w58_0_c0 & bh59_w57_0_c0 & bh59_w56_0_c0 & bh59_w55_0_c0 & bh59_w54_0_c0 & bh59_w53_0_c0 & bh59_w52_0_c0 & bh59_w51_0_c0 & bh59_w50_0_c0 & bh59_w49_0_c0 & bh59_w48_0_c0 & bh59_w47_0_c0 & bh59_w46_0_c0 & bh59_w45_0_c0 & bh59_w44_0_c0 & bh59_w43_0_c0 & bh59_w42_0_c0 & bh59_w41_0_c0 & bh59_w40_0_c0 & bh59_w39_0_c0 & bh59_w38_0_c0 & bh59_w37_0_c0 & bh59_w36_0_c0 & bh59_w35_0_c0 & bh59_w34_0_c0 & bh59_w33_0_c0 & bh59_w32_0_c0 & bh59_w31_0_c0 & bh59_w30_0_c0 & bh59_w29_0_c0 & bh59_w28_0_c0 & bh59_w27_0_c0 & bh59_w26_0_c0 & bh59_w25_0_c0 & bh59_w24_0_c0 & bh59_w23_0_c0 & bh59_w22_0_c0 & bh59_w21_0_c0 & bh59_w20_0_c0 & bh59_w19_0_c0 & bh59_w18_0_c0 & bh59_w17_0_c0 & bh59_w16_0_c0 & bh59_w15_0_c0 & bh59_w14_0_c0 & bh59_w13_0_c0 & bh59_w12_0_c0 & bh59_w11_0_c0 & bh59_w10_0_c0 & bh59_w9_0_c0 & bh59_w8_0_c0 & bh59_w7_0_c0 & bh59_w6_0_c0 & bh59_w5_0_c0 & bh59_w4_0_c0 & bh59_w3_0_c0 & bh59_w2_0_c0 & bh59_w1_0_c0 & bh59_w0_0_c0;
   bitheapFinalAdd_bh59_In1_c0 <= "0" & "0" & "0" & "0" & "0" & "0" & bh59_w75_1_c0 & bh59_w74_1_c0 & bh59_w73_1_c0 & bh59_w72_1_c0 & bh59_w71_1_c0 & bh59_w70_1_c0 & bh59_w69_1_c0 & bh59_w68_1_c0 & bh59_w67_1_c0 & bh59_w66_1_c0 & bh59_w65_1_c0 & bh59_w64_1_c0 & bh59_w63_1_c0 & bh59_w62_1_c0 & bh59_w61_1_c0 & bh59_w60_1_c0 & bh59_w59_1_c0 & bh59_w58_1_c0 & bh59_w57_1_c0 & bh59_w56_1_c0 & bh59_w55_1_c0 & bh59_w54_1_c0 & bh59_w53_1_c0 & bh59_w52_1_c0 & bh59_w51_1_c0 & bh59_w50_1_c0 & bh59_w49_1_c0 & bh59_w48_1_c0 & bh59_w47_1_c0 & bh59_w46_1_c0 & bh59_w45_1_c0 & bh59_w44_1_c0 & bh59_w43_1_c0 & bh59_w42_1_c0 & bh59_w41_1_c0 & bh59_w40_1_c0 & bh59_w39_1_c0 & bh59_w38_1_c0 & bh59_w37_1_c0 & bh59_w36_1_c0 & bh59_w35_1_c0 & bh59_w34_1_c0 & bh59_w33_1_c0 & bh59_w32_1_c0 & bh59_w31_1_c0 & bh59_w30_1_c0 & bh59_w29_1_c0 & bh59_w28_1_c0 & bh59_w27_1_c0 & bh59_w26_1_c0 & bh59_w25_1_c0 & bh59_w24_1_c0 & bh59_w23_1_c0 & bh59_w22_1_c0 & bh59_w21_1_c0 & bh59_w20_1_c0 & bh59_w19_1_c0 & bh59_w18_1_c0 & bh59_w17_1_c0 & bh59_w16_1_c0 & bh59_w15_1_c0 & bh59_w14_1_c0 & bh59_w13_1_c0 & bh59_w12_1_c0 & bh59_w11_1_c0 & bh59_w10_1_c0 & bh59_w9_1_c0 & bh59_w8_1_c0 & bh59_w7_1_c0 & bh59_w6_1_c0 & bh59_w5_1_c0 & bh59_w4_1_c0 & bh59_w3_1_c0 & bh59_w2_1_c0 & bh59_w1_1_c0 & bh59_w0_1_c0;
   bitheapFinalAdd_bh59_Cin_c0 <= '0';

   bitheapFinalAdd_bh59: IntAdder_82_Freq300_uid68
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 Cin => bitheapFinalAdd_bh59_Cin_c0,
                 X => bitheapFinalAdd_bh59_In0_c0,
                 Y => bitheapFinalAdd_bh59_In1_c0,
                 R => bitheapFinalAdd_bh59_Out_c1);
   bitheapResult_bh59_c1 <= bitheapFinalAdd_bh59_Out_c1(80 downto 0);
   OutRes_c1 <= bitheapResult_bh59_c1(80 downto 0);
   R <= OutRes_c1(80 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_115_Freq300_uid70
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_115_Freq300_uid70 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(114 downto 0);
          Y : in  std_logic_vector(114 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(114 downto 0)   );
end entity;

architecture arch of IntAdder_115_Freq300_uid70 is
signal Rtmp_c9 :  std_logic_vector(114 downto 0);
signal X_c2, X_c3, X_c4, X_c5, X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(114 downto 0);
signal Y_c9 :  std_logic_vector(114 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               X_c2 <= X;
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               X_c3 <= X_c2;
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               X_c4 <= X_c3;
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               X_c5 <= X_c4;
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
               Y_c9 <= Y;
               Cin_c9 <= Cin_c8;
            end if;
         end if;
      end process;
   Rtmp_c9 <= X_c9 + Y_c9 + Cin_c9;
   R <= Rtmp_c9;
end architecture;

--------------------------------------------------------------------------------
--                   Normalizer_Z_115_104_44_Freq300_uid72
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_115_104_44_Freq300_uid72 is
    port (clk, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(114 downto 0);
          Count : out  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(103 downto 0)   );
end entity;

architecture arch of Normalizer_Z_115_104_44_Freq300_uid72 is
signal level6_c9 :  std_logic_vector(114 downto 0);
signal count5_c9, count5_c10, count5_c11 :  std_logic;
signal level5_c9 :  std_logic_vector(114 downto 0);
signal count4_c9, count4_c10, count4_c11 :  std_logic;
signal level4_c9, level4_c10 :  std_logic_vector(114 downto 0);
signal count3_c9, count3_c10, count3_c11 :  std_logic;
signal level3_c10 :  std_logic_vector(110 downto 0);
signal count2_c10, count2_c11 :  std_logic;
signal level2_c10 :  std_logic_vector(106 downto 0);
signal count1_c10, count1_c11 :  std_logic;
signal level1_c10, level1_c11 :  std_logic_vector(104 downto 0);
signal count0_c11 :  std_logic;
signal level0_c11 :  std_logic_vector(103 downto 0);
signal sCount_c11 :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_10 = '1' then
               count5_c10 <= count5_c9;
               count4_c10 <= count4_c9;
               level4_c10 <= level4_c9;
               count3_c10 <= count3_c9;
            end if;
            if ce_11 = '1' then
               count5_c11 <= count5_c10;
               count4_c11 <= count4_c10;
               count3_c11 <= count3_c10;
               count2_c11 <= count2_c10;
               count1_c11 <= count1_c10;
               level1_c11 <= level1_c10;
            end if;
         end if;
      end process;
   level6_c9 <= X ;
   count5_c9<= '1' when level6_c9(114 downto 83) = (114 downto 83=>'0') else '0';
   level5_c9<= level6_c9(114 downto 0) when count5_c9='0' else level6_c9(82 downto 0) & (31 downto 0 => '0');

   count4_c9<= '1' when level5_c9(114 downto 99) = (114 downto 99=>'0') else '0';
   level4_c9<= level5_c9(114 downto 0) when count4_c9='0' else level5_c9(98 downto 0) & (15 downto 0 => '0');

   count3_c9<= '1' when level4_c9(114 downto 107) = (114 downto 107=>'0') else '0';
   level3_c10<= level4_c10(114 downto 4) when count3_c10='0' else level4_c10(106 downto 0) & (3 downto 0 => '0');

   count2_c10<= '1' when level3_c10(110 downto 107) = (110 downto 107=>'0') else '0';
   level2_c10<= level3_c10(110 downto 4) when count2_c10='0' else level3_c10(106 downto 0);

   count1_c10<= '1' when level2_c10(106 downto 105) = (106 downto 105=>'0') else '0';
   level1_c10<= level2_c10(106 downto 2) when count1_c10='0' else level2_c10(104 downto 0);

   count0_c11<= '1' when level1_c11(104 downto 104) = (104 downto 104=>'0') else '0';
   level0_c11<= level1_c11(104 downto 1) when count0_c11='0' else level1_c11(103 downto 0);

   R <= level0_c11;
   sCount_c11 <= count5_c11 & count4_c11 & count3_c11 & count2_c11 & count1_c11 & count0_c11;
   Count <= sCount_c11;
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter38_by_max_37_Freq300_uid74
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X S
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter38_by_max_37_Freq300_uid74 is
    port (clk, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(37 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(74 downto 0)   );
end entity;

architecture arch of RightShifter38_by_max_37_Freq300_uid74 is
signal ps_c3, ps_c4, ps_c5, ps_c6, ps_c7, ps_c8 :  std_logic_vector(5 downto 0);
signal level0_c6 :  std_logic_vector(37 downto 0);
signal level1_c6, level1_c7 :  std_logic_vector(38 downto 0);
signal level2_c7 :  std_logic_vector(40 downto 0);
signal level3_c7 :  std_logic_vector(44 downto 0);
signal level4_c7 :  std_logic_vector(52 downto 0);
signal level5_c7, level5_c8 :  std_logic_vector(68 downto 0);
signal level6_c8 :  std_logic_vector(100 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_4 = '1' then
               ps_c4 <= ps_c3;
            end if;
            if ce_5 = '1' then
               ps_c5 <= ps_c4;
            end if;
            if ce_6 = '1' then
               ps_c6 <= ps_c5;
            end if;
            if ce_7 = '1' then
               ps_c7 <= ps_c6;
               level1_c7 <= level1_c6;
            end if;
            if ce_8 = '1' then
               ps_c8 <= ps_c7;
               level5_c8 <= level5_c7;
            end if;
         end if;
      end process;
   ps_c3<= S;
   level0_c6<= X;
   level1_c6 <=  (0 downto 0 => '0') & level0_c6 when ps_c6(0) = '1' else    level0_c6 & (0 downto 0 => '0');
   level2_c7 <=  (1 downto 0 => '0') & level1_c7 when ps_c7(1) = '1' else    level1_c7 & (1 downto 0 => '0');
   level3_c7 <=  (3 downto 0 => '0') & level2_c7 when ps_c7(2) = '1' else    level2_c7 & (3 downto 0 => '0');
   level4_c7 <=  (7 downto 0 => '0') & level3_c7 when ps_c7(3) = '1' else    level3_c7 & (7 downto 0 => '0');
   level5_c7 <=  (15 downto 0 => '0') & level4_c7 when ps_c7(4) = '1' else    level4_c7 & (15 downto 0 => '0');
   level6_c8 <=  (31 downto 0 => '0') & level5_c8 when ps_c8(5) = '1' else    level5_c8 & (31 downto 0 => '0');
   R <= level6_c8(100 downto 26);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_72_Freq300_uid76
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_72_Freq300_uid76 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(71 downto 0);
          Y : in  std_logic_vector(71 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(71 downto 0)   );
end entity;

architecture arch of IntAdder_72_Freq300_uid76 is
signal Rtmp_c8 :  std_logic_vector(71 downto 0);
signal X_c5, X_c6, X_c7, X_c8 :  std_logic_vector(71 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               X_c5 <= X;
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
               Cin_c8 <= Cin_c7;
            end if;
         end if;
      end process;
   Rtmp_c8 <= X_c8 + Y + Cin_c8;
   R <= Rtmp_c8;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_77_Freq300_uid79
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_77_Freq300_uid79 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(76 downto 0);
          Y : in  std_logic_vector(76 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(76 downto 0)   );
end entity;

architecture arch of IntAdder_77_Freq300_uid79 is
signal Rtmp_c11 :  std_logic_vector(76 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
         end if;
      end process;
   Rtmp_c11 <= X + Y + Cin_c11;
   R <= Rtmp_c11;
end architecture;

--------------------------------------------------------------------------------
--                  FPLogIterative_11_66_0_300_Freq300_uid9
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPLogIterative_11_66_0_300_Freq300_uid9 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(11+66+2 downto 0);
          R : out  std_logic_vector(11+66+2 downto 0)   );
end entity;

architecture arch of FPLogIterative_11_66_0_300_Freq300_uid9 is
   component LZOC_66_Freq300_uid11 is
      port ( clk, ce_1, ce_2 : in std_logic;
             I : in  std_logic_vector(65 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(6 downto 0)   );
   end component;

   component LeftShifter34_by_max_34_Freq300_uid13 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(33 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(67 downto 0)   );
   end component;

   component InvA0Table_Freq300_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component IntAdder_80_Freq300_uid18 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(79 downto 0);
             Y : in  std_logic_vector(79 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(79 downto 0)   );
   end component;

   component IntAdder_80_Freq300_uid21 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(79 downto 0);
             Y : in  std_logic_vector(79 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(79 downto 0)   );
   end component;

   component IntAdder_79_Freq300_uid24 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(78 downto 0);
             Y : in  std_logic_vector(78 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(78 downto 0)   );
   end component;

   component IntAdder_79_Freq300_uid27 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(78 downto 0);
             Y : in  std_logic_vector(78 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(78 downto 0)   );
   end component;

   component IntAdder_70_Freq300_uid30 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(69 downto 0);
             Y : in  std_logic_vector(69 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(69 downto 0)   );
   end component;

   component IntAdder_70_Freq300_uid33 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(69 downto 0);
             Y : in  std_logic_vector(69 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(69 downto 0)   );
   end component;

   component IntAdder_70_Freq300_uid36 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7 : in std_logic;
             X : in  std_logic_vector(69 downto 0);
             Y : in  std_logic_vector(69 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(69 downto 0)   );
   end component;

   component LogTable0_Freq300_uid38 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : out  std_logic_vector(103 downto 0)   );
   end component;

   component LogTable1_Freq300_uid40 is
      port ( clk, ce_2 : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(94 downto 0)   );
   end component;

   component IntAdder_104_Freq300_uid43 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(103 downto 0);
             Y : in  std_logic_vector(103 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(103 downto 0)   );
   end component;

   component LogTable2_Freq300_uid45 is
      port ( clk, ce_4 : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(86 downto 0)   );
   end component;

   component IntAdder_104_Freq300_uid48 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(103 downto 0);
             Y : in  std_logic_vector(103 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(103 downto 0)   );
   end component;

   component LogTable3_Freq300_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(78 downto 0)   );
   end component;

   component IntAdder_104_Freq300_uid53 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(103 downto 0);
             Y : in  std_logic_vector(103 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(103 downto 0)   );
   end component;

   component IntAdder_104_Freq300_uid56 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(103 downto 0);
             Y : in  std_logic_vector(103 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(103 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid58 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             R : out  std_logic_vector(80 downto 0)   );
   end component;

   component IntAdder_115_Freq300_uid70 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(114 downto 0);
             Y : in  std_logic_vector(114 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(114 downto 0)   );
   end component;

   component Normalizer_Z_115_104_44_Freq300_uid72 is
      port ( clk, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(114 downto 0);
             Count : out  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(103 downto 0)   );
   end component;

   component RightShifter38_by_max_37_Freq300_uid74 is
      port ( clk, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(37 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(74 downto 0)   );
   end component;

   component IntAdder_72_Freq300_uid76 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(71 downto 0);
             Y : in  std_logic_vector(71 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(71 downto 0)   );
   end component;

   component IntAdder_77_Freq300_uid79 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(76 downto 0);
             Y : in  std_logic_vector(76 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(76 downto 0)   );
   end component;

signal XExnSgn_c0, XExnSgn_c1, XExnSgn_c2, XExnSgn_c3, XExnSgn_c4, XExnSgn_c5, XExnSgn_c6, XExnSgn_c7, XExnSgn_c8, XExnSgn_c9, XExnSgn_c10, XExnSgn_c11 :  std_logic_vector(2 downto 0);
signal FirstBit_c0 :  std_logic;
signal Y0_c0, Y0_c1 :  std_logic_vector(67 downto 0);
signal Y0h_c0 :  std_logic_vector(65 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6, sR_c7, sR_c8, sR_c9, sR_c10, sR_c11 :  std_logic;
signal absZ0_c0 :  std_logic_vector(33 downto 0);
signal E_c0 :  std_logic_vector(10 downto 0);
signal absE_c0 :  std_logic_vector(10 downto 0);
signal EeqZero_c0, EeqZero_c1, EeqZero_c2, EeqZero_c3 :  std_logic;
signal lzo_c2, lzo_c3, lzo_c4, lzo_c5, lzo_c6, lzo_c7, lzo_c8 :  std_logic_vector(6 downto 0);
signal pfinal_s_c0, pfinal_s_c1, pfinal_s_c2, pfinal_s_c3 :  std_logic_vector(6 downto 0);
signal shiftval_c3 :  std_logic_vector(7 downto 0);
signal shiftvalinL_c3 :  std_logic_vector(5 downto 0);
signal shiftvalinR_c3 :  std_logic_vector(5 downto 0);
signal doRR_c3, doRR_c4, doRR_c5, doRR_c6 :  std_logic;
signal small_c3, small_c4, small_c5, small_c6, small_c7, small_c8, small_c9, small_c10, small_c11 :  std_logic;
signal small_absZ0_normd_full_c4 :  std_logic_vector(67 downto 0);
signal small_absZ0_normd_c4, small_absZ0_normd_c5, small_absZ0_normd_c6 :  std_logic_vector(33 downto 0);
signal A0_c0 :  std_logic_vector(10 downto 0);
signal InvA0_c0, InvA0_c1 :  std_logic_vector(11 downto 0);
signal P0_c1 :  std_logic_vector(79 downto 0);
signal Z1_c1 :  std_logic_vector(68 downto 0);
signal A1_c1, A1_c2 :  std_logic_vector(8 downto 0);
signal B1_c1 :  std_logic_vector(59 downto 0);
signal ZM1_c1, ZM1_c2 :  std_logic_vector(68 downto 0);
signal P1_c2 :  std_logic_vector(77 downto 0);
signal Y1_c1 :  std_logic_vector(78 downto 0);
signal EiY1_c1 :  std_logic_vector(79 downto 0);
signal addXIter1_c1 :  std_logic_vector(79 downto 0);
signal EiYPB1_c2 :  std_logic_vector(79 downto 0);
signal Pp1_c2 :  std_logic_vector(79 downto 0);
signal Z2_c3 :  std_logic_vector(79 downto 0);
signal A2_c3, A2_c4 :  std_logic_vector(8 downto 0);
signal B2_c3 :  std_logic_vector(70 downto 0);
signal ZM2_c3, ZM2_c4 :  std_logic_vector(69 downto 0);
signal P2_c4 :  std_logic_vector(78 downto 0);
signal Y2_c3 :  std_logic_vector(97 downto 0);
signal EiY2_c3 :  std_logic_vector(78 downto 0);
signal addXIter2_c3 :  std_logic_vector(78 downto 0);
signal EiYPB2_c4 :  std_logic_vector(78 downto 0);
signal Pp2_c4 :  std_logic_vector(78 downto 0);
signal Z3_c5 :  std_logic_vector(78 downto 0);
signal A3_c5 :  std_logic_vector(9 downto 0);
signal B3_c5 :  std_logic_vector(68 downto 0);
signal ZM3_c5 :  std_logic_vector(53 downto 0);
signal P3_c5, P3_c6 :  std_logic_vector(63 downto 0);
signal Y3_c5 :  std_logic_vector(104 downto 0);
signal EiY3_c5 :  std_logic_vector(69 downto 0);
signal addXIter3_c5 :  std_logic_vector(69 downto 0);
signal EiYPB3_c5 :  std_logic_vector(69 downto 0);
signal Pp3_c6 :  std_logic_vector(69 downto 0);
signal Z4_c6 :  std_logic_vector(69 downto 0);
signal Zfinal_c6 :  std_logic_vector(69 downto 0);
signal squarerIn_c6 :  std_logic_vector(37 downto 0);
signal Z2o2_full_c6 :  std_logic_vector(75 downto 0);
signal Z2o2_full_dummy_c6 :  std_logic_vector(75 downto 0);
signal Z2o2_normal_c6 :  std_logic_vector(34 downto 0);
signal addFinalLog1pY_c6 :  std_logic_vector(69 downto 0);
signal Log1p_normal_c7 :  std_logic_vector(69 downto 0);
signal L0_c0 :  std_logic_vector(103 downto 0);
signal S1_c0 :  std_logic_vector(103 downto 0);
signal L1_c2 :  std_logic_vector(94 downto 0);
signal sopX1_c2 :  std_logic_vector(103 downto 0);
signal S2_c2 :  std_logic_vector(103 downto 0);
signal L2_c4 :  std_logic_vector(86 downto 0);
signal sopX2_c4 :  std_logic_vector(103 downto 0);
signal S3_c4 :  std_logic_vector(103 downto 0);
signal L3_c5 :  std_logic_vector(78 downto 0);
signal sopX3_c5 :  std_logic_vector(103 downto 0);
signal S4_c6 :  std_logic_vector(103 downto 0);
signal almostLog_c6 :  std_logic_vector(103 downto 0);
signal adderLogF_normalY_c7 :  std_logic_vector(103 downto 0);
signal LogF_normal_c8 :  std_logic_vector(103 downto 0);
signal absELog2_c1 :  std_logic_vector(80 downto 0);
signal absELog2_pad_c1 :  std_logic_vector(114 downto 0);
signal LogF_normal_pad_c8 :  std_logic_vector(114 downto 0);
signal lnaddX_c1 :  std_logic_vector(114 downto 0);
signal lnaddY_c8 :  std_logic_vector(114 downto 0);
signal Log_normal_c9 :  std_logic_vector(114 downto 0);
signal Log_normal_normd_c11 :  std_logic_vector(103 downto 0);
signal E_normal_c11 :  std_logic_vector(5 downto 0);
signal Z2o2_small_bs_c6 :  std_logic_vector(37 downto 0);
signal Z2o2_small_s_c8 :  std_logic_vector(74 downto 0);
signal Z2o2_small_c8 :  std_logic_vector(71 downto 0);
signal Z_small_c4 :  std_logic_vector(71 downto 0);
signal Log_smallY_c8 :  std_logic_vector(71 downto 0);
signal nsRCin_c0 :  std_logic;
signal Log_small_c8 :  std_logic_vector(71 downto 0);
signal E0_sub_c8 :  std_logic_vector(1 downto 0);
signal ufl_c0, ufl_c1, ufl_c2, ufl_c3, ufl_c4, ufl_c5, ufl_c6, ufl_c7, ufl_c8, ufl_c9, ufl_c10, ufl_c11 :  std_logic;
signal E_small_c8, E_small_c9, E_small_c10, E_small_c11 :  std_logic_vector(10 downto 0);
signal Log_small_normd_c8, Log_small_normd_c9, Log_small_normd_c10, Log_small_normd_c11 :  std_logic_vector(69 downto 0);
signal E0offset_c0, E0offset_c1, E0offset_c2, E0offset_c3, E0offset_c4, E0offset_c5, E0offset_c6, E0offset_c7, E0offset_c8, E0offset_c9, E0offset_c10, E0offset_c11 :  std_logic_vector(10 downto 0);
signal ER_c11 :  std_logic_vector(10 downto 0);
signal Log_g_c11 :  std_logic_vector(69 downto 0);
signal round_c11 :  std_logic;
signal fraX_c11 :  std_logic_vector(76 downto 0);
signal fraY_c11 :  std_logic_vector(76 downto 0);
signal EFR_c11 :  std_logic_vector(76 downto 0);
signal Rexn_c11 :  std_logic_vector(2 downto 0);
constant g: positive := 4;
constant log2wF: positive := 7;
constant pfinal: positive := 34;
constant sfinal: positive := 70;
constant targetprec: positive := 104;
constant wE: positive := 11;
constant wF: positive := 66;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               XExnSgn_c1 <= XExnSgn_c0;
               Y0_c1 <= Y0_c0;
               sR_c1 <= sR_c0;
               EeqZero_c1 <= EeqZero_c0;
               pfinal_s_c1 <= pfinal_s_c0;
               InvA0_c1 <= InvA0_c0;
               ufl_c1 <= ufl_c0;
               E0offset_c1 <= E0offset_c0;
            end if;
            if ce_2 = '1' then
               XExnSgn_c2 <= XExnSgn_c1;
               sR_c2 <= sR_c1;
               EeqZero_c2 <= EeqZero_c1;
               pfinal_s_c2 <= pfinal_s_c1;
               A1_c2 <= A1_c1;
               ZM1_c2 <= ZM1_c1;
               ufl_c2 <= ufl_c1;
               E0offset_c2 <= E0offset_c1;
            end if;
            if ce_3 = '1' then
               XExnSgn_c3 <= XExnSgn_c2;
               sR_c3 <= sR_c2;
               EeqZero_c3 <= EeqZero_c2;
               lzo_c3 <= lzo_c2;
               pfinal_s_c3 <= pfinal_s_c2;
               ufl_c3 <= ufl_c2;
               E0offset_c3 <= E0offset_c2;
            end if;
            if ce_4 = '1' then
               XExnSgn_c4 <= XExnSgn_c3;
               sR_c4 <= sR_c3;
               lzo_c4 <= lzo_c3;
               doRR_c4 <= doRR_c3;
               small_c4 <= small_c3;
               A2_c4 <= A2_c3;
               ZM2_c4 <= ZM2_c3;
               ufl_c4 <= ufl_c3;
               E0offset_c4 <= E0offset_c3;
            end if;
            if ce_5 = '1' then
               XExnSgn_c5 <= XExnSgn_c4;
               sR_c5 <= sR_c4;
               lzo_c5 <= lzo_c4;
               doRR_c5 <= doRR_c4;
               small_c5 <= small_c4;
               small_absZ0_normd_c5 <= small_absZ0_normd_c4;
               ufl_c5 <= ufl_c4;
               E0offset_c5 <= E0offset_c4;
            end if;
            if ce_6 = '1' then
               XExnSgn_c6 <= XExnSgn_c5;
               sR_c6 <= sR_c5;
               lzo_c6 <= lzo_c5;
               doRR_c6 <= doRR_c5;
               small_c6 <= small_c5;
               small_absZ0_normd_c6 <= small_absZ0_normd_c5;
               P3_c6 <= P3_c5;
               ufl_c6 <= ufl_c5;
               E0offset_c6 <= E0offset_c5;
            end if;
            if ce_7 = '1' then
               XExnSgn_c7 <= XExnSgn_c6;
               sR_c7 <= sR_c6;
               lzo_c7 <= lzo_c6;
               small_c7 <= small_c6;
               ufl_c7 <= ufl_c6;
               E0offset_c7 <= E0offset_c6;
            end if;
            if ce_8 = '1' then
               XExnSgn_c8 <= XExnSgn_c7;
               sR_c8 <= sR_c7;
               lzo_c8 <= lzo_c7;
               small_c8 <= small_c7;
               ufl_c8 <= ufl_c7;
               E0offset_c8 <= E0offset_c7;
            end if;
            if ce_9 = '1' then
               XExnSgn_c9 <= XExnSgn_c8;
               sR_c9 <= sR_c8;
               small_c9 <= small_c8;
               ufl_c9 <= ufl_c8;
               E_small_c9 <= E_small_c8;
               Log_small_normd_c9 <= Log_small_normd_c8;
               E0offset_c9 <= E0offset_c8;
            end if;
            if ce_10 = '1' then
               XExnSgn_c10 <= XExnSgn_c9;
               sR_c10 <= sR_c9;
               small_c10 <= small_c9;
               ufl_c10 <= ufl_c9;
               E_small_c10 <= E_small_c9;
               Log_small_normd_c10 <= Log_small_normd_c9;
               E0offset_c10 <= E0offset_c9;
            end if;
            if ce_11 = '1' then
               XExnSgn_c11 <= XExnSgn_c10;
               sR_c11 <= sR_c10;
               small_c11 <= small_c10;
               ufl_c11 <= ufl_c10;
               E_small_c11 <= E_small_c10;
               Log_small_normd_c11 <= Log_small_normd_c10;
               E0offset_c11 <= E0offset_c10;
            end if;
         end if;
      end process;
   XExnSgn_c0 <=  X(wE+wF+2 downto wE+wF);
   FirstBit_c0 <=  X(wF-1);
   Y0_c0 <= "1" & X(wF-1 downto 0) & "0" when FirstBit_c0 = '0' else "01" & X(wF-1 downto 0);
   Y0h_c0 <= Y0_c0(wF downto 1);
   -- Sign of the result;
   sR_c0 <= '0'   when  (X(wE+wF-1 downto wF) = ('0' & (wE-2 downto 0 => '1')))  -- binade [1..2)
     else not X(wE+wF-1);                -- MSB of exponent
   absZ0_c0 <=   Y0_c0(wF-pfinal+1 downto 0)          when (sR_c0='0') else
             ((wF-pfinal+1 downto 0 => '0') - Y0_c0(wF-pfinal+1 downto 0));
   E_c0 <= (X(wE+wF-1 downto wF)) - ("0" & (wE-2 downto 1 => '1') & (not FirstBit_c0));
   absE_c0 <= ((wE-1 downto 0 => '0') - E_c0)   when sR_c0 = '1' else E_c0;
   EeqZero_c0 <= '1' when E_c0=(wE-1 downto 0 => '0') else '0';
   lzoc1: LZOC_66_Freq300_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 I => Y0h_c0,
                 OZB => FirstBit_c0,
                 O => lzo_c2);
   pfinal_s_c0 <= "0100010";
   shiftval_c3 <= ('0' & lzo_c3) - ('0' & pfinal_s_c3); 
   shiftvalinL_c3 <= shiftval_c3(5 downto 0);
   shiftvalinR_c3 <= shiftval_c3(5 downto 0);
   doRR_c3 <= shiftval_c3(log2wF); -- sign of the result
   small_c3 <= EeqZero_c3 and not(doRR_c3);
   -- The left shifter for the 'small' case
   small_lshift: LeftShifter34_by_max_34_Freq300_uid13
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 S => shiftvalinL_c3,
                 X => absZ0_c0,
                 R => small_absZ0_normd_full_c4);
   small_absZ0_normd_c4 <= small_absZ0_normd_full_c4(33 downto 0); -- get rid of leading zeroes
   ---------------- The range reduction box ---------------
   A0_c0 <= X(65 downto 55);
   -- First inv table
   InvA0Table: InvA0Table_Freq300_uid15
      port map ( clk  => clk,
                 X => A0_c0,
                 Y => InvA0_c0);
   P0_c1 <= InvA0_c1 * Y0_c1;

   Z1_c1 <= P0_c1(68 downto 0);

   A1_c1 <= Z1_c1(68 downto 60);
   B1_c1 <= Z1_c1(59 downto 0);
   ZM1_c1 <= Z1_c1;
   P1_c2 <= A1_c2*ZM1_c2;
   Y1_c1 <= "1" & (8 downto 0 => '0') & Z1_c1;
   EiY1_c1 <= Y1_c1 & (0 downto 0 => '0')  when A1_c1(8) = '1'
     else  "0" & Y1_c1;
   addXIter1_c1 <= "0" & B1_c1 & (18 downto 0 => '0');
   addIter1_1: IntAdder_80_Freq300_uid18
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => '0',
                 X => addXIter1_c1,
                 Y => EiY1_c1,
                 R => EiYPB1_c2);
   Pp1_c2 <= (0 downto 0 => '1') & not(P1_c2 & (0 downto 0 => '0'));
   addIter2_1: IntAdder_80_Freq300_uid21
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 Cin => '1',
                 X => EiYPB1_c2,
                 Y => Pp1_c2,
                 R => Z2_c3);

   A2_c3 <= Z2_c3(79 downto 71);
   B2_c3 <= Z2_c3(70 downto 0);
   ZM2_c3 <= Z2_c3(79 downto 10);
   P2_c4 <= A2_c4*ZM2_c4;
   Y2_c3 <= "1" & (16 downto 0 => '0') & Z2_c3;
   EiY2_c3 <= (7 downto 0 => '0') & Y2_c3(97 downto 27);
   addXIter2_c3 <= "0" & B2_c3 & (6 downto 0 => '0');
   addIter1_2: IntAdder_79_Freq300_uid24
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 Cin => '0',
                 X => addXIter2_c3,
                 Y => EiY2_c3,
                 R => EiYPB2_c4);
   Pp2_c4 <= (8 downto 0 => '1') & not(P2_c4(78 downto 9));
   addIter2_2: IntAdder_79_Freq300_uid27
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 Cin => '1',
                 X => EiYPB2_c4,
                 Y => Pp2_c4,
                 R => Z3_c5);

   A3_c5 <= Z3_c5(78 downto 69);
   B3_c5 <= Z3_c5(68 downto 0);
   ZM3_c5 <= Z3_c5(78 downto 25);
   P3_c5 <= A3_c5*ZM3_c5;
   Y3_c5 <= "1" & (24 downto 0 => '0') & Z3_c5;
   EiY3_c5 <= (14 downto 0 => '0') & Y3_c5(104 downto 50);
   addXIter3_c5 <= "0" & B3_c5;
   addIter1_3: IntAdder_70_Freq300_uid30
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 Cin => '0',
                 X => addXIter3_c5,
                 Y => EiY3_c5,
                 R => EiYPB3_c5);
   Pp3_c6 <= (15 downto 0 => '1') & not(P3_c6(63 downto 10));
   addIter2_3: IntAdder_70_Freq300_uid33
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 Cin => '1',
                 X => EiYPB3_c5,
                 Y => Pp3_c6,
                 R => Z4_c6);
   Zfinal_c6 <= Z4_c6;
   squarerIn_c6 <= Zfinal_c6(sfinal-1 downto sfinal-38) when doRR_c6='1'
                    else (small_absZ0_normd_c6 & (3 downto 0 => '0'));  
   Z2o2_full_c6 <= squarerIn_c6*squarerIn_c6;
   Z2o2_full_dummy_c6 <= Z2o2_full_c6;
   Z2o2_normal_c6 <= Z2o2_full_dummy_c6 (75  downto 41);
   addFinalLog1pY_c6 <= (pfinal downto 0  => '1') & not(Z2o2_normal_c6);
   addFinalLog1p_normalAdder: IntAdder_70_Freq300_uid36
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 Cin => '1',
                 X => Zfinal_c6,
                 Y => addFinalLog1pY_c6,
                 R => Log1p_normal_c7);

   -- Now the log tables, as late as possible
   LogTable0: LogTable0_Freq300_uid38
      port map ( clk  => clk,
                 X => A0_c0,
                 Y => L0_c0);
   S1_c0 <= L0_c0;
   LogTable1: LogTable1_Freq300_uid40
      port map ( clk  => clk,
                 ce_2 => ce_2,
                 X => A1_c1,
                 Y => L1_c2);
   sopX1_c2 <= ((103 downto 95 => '0') & L1_c2);
   adderS1: IntAdder_104_Freq300_uid43
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => '0',
                 X => S1_c0,
                 Y => sopX1_c2,
                 R => S2_c2);
   LogTable2: LogTable2_Freq300_uid45
      port map ( clk  => clk,
                 ce_4 => ce_4,
                 X => A2_c3,
                 Y => L2_c4);
   sopX2_c4 <= ((103 downto 87 => '0') & L2_c4);
   adderS2: IntAdder_104_Freq300_uid48
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 Cin => '0',
                 X => S2_c2,
                 Y => sopX2_c4,
                 R => S3_c4);
   LogTable3: LogTable3_Freq300_uid50
      port map ( clk  => clk,
                 X => A3_c5,
                 Y => L3_c5);
   sopX3_c5 <= ((103 downto 79 => '0') & L3_c5);
   adderS3: IntAdder_104_Freq300_uid53
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 Cin => '0',
                 X => S3_c4,
                 Y => sopX3_c5,
                 R => S4_c6);
   almostLog_c6 <= S4_c6;
   adderLogF_normalY_c7 <= ((targetprec-1 downto sfinal => '0') & Log1p_normal_c7);
   adderLogF_normal: IntAdder_104_Freq300_uid56
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 Cin => '0',
                 X => almostLog_c6,
                 Y => adderLogF_normalY_c7,
                 R => LogF_normal_c8);
   MulLog2: FixRealKCM_Freq300_uid58
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => absE_c0,
                 R => absELog2_c1);
   absELog2_pad_c1 <=   absELog2_c1 & (targetprec-wF-g-1 downto 0 => '0');       
   LogF_normal_pad_c8 <= (wE-1  downto 0 => LogF_normal_c8(targetprec-1))  & LogF_normal_c8;
   lnaddX_c1 <= absELog2_pad_c1;
   lnaddY_c8 <= LogF_normal_pad_c8 when sR_c8='0' else not(LogF_normal_pad_c8); 
   lnadder: IntAdder_115_Freq300_uid70
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 Cin => sR_c0,
                 X => lnaddX_c1,
                 Y => lnaddY_c8,
                 R => Log_normal_c9);
   final_norm: Normalizer_Z_115_104_44_Freq300_uid72
      port map ( clk  => clk,
                 ce_10 => ce_10,
                 ce_11=> ce_11,
                 X => Log_normal_c9,
                 Count => E_normal_c11,
                 R => Log_normal_normd_c11);
   Z2o2_small_bs_c6 <= Z2o2_full_dummy_c6(75 downto 38);
   ao_rshift: RightShifter38_by_max_37_Freq300_uid74
      port map ( clk  => clk,
                 ce_4 => ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 S => shiftvalinR_c3,
                 X => Z2o2_small_bs_c6,
                 R => Z2o2_small_s_c8);
     -- send the MSB to position pfinal
   Z2o2_small_c8 <=  (pfinal-1 downto 0  => '0') & Z2o2_small_s_c8(74 downto 37);
   -- mantissa will be either Y0-z^2/2  or  -Y0+z^2/2,  depending on sR  
   Z_small_c4 <= small_absZ0_normd_c4 & (37 downto 0 => '0');
   Log_smallY_c8 <= Z2o2_small_c8 when sR_c8='1' else not(Z2o2_small_c8);
   nsRCin_c0 <= not ( sR_c0 );
   log_small_adder: IntAdder_72_Freq300_uid76
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 Cin => nsRCin_c0,
                 X => Z_small_c4,
                 Y => Log_smallY_c8,
                 R => Log_small_c8);
   -- Possibly subtract 1 or 2 to the exponent, depending on the LZC of Log_small
   E0_sub_c8 <=   "11" when Log_small_c8(wF+g+1) = '1'
          else "10" when Log_small_c8(wF+g+1 downto wF+g) = "01"
          else "01" ;
   -- The smallest log will be log(1+2^{-wF}) \approx 2^{-wF}  = 2^-66
   -- The smallest representable number is 2^{1-2^(wE-1)} = 2^-1023
   -- No underflow possible
   ufl_c0 <= '0';
   E_small_c8 <=  ("0" & (wE-2 downto 2 => '1') & E0_sub_c8)  -  ((wE-1 downto 7 => '0') & lzo_c8) ;
   Log_small_normd_c8 <= Log_small_c8(wF+g+1 downto 2) when Log_small_c8(wF+g+1)='1'
           else Log_small_c8(wF+g downto 1)  when Log_small_c8(wF+g)='1'  -- remove the first zero
           else Log_small_c8(wF+g-1 downto 0)  ; -- remove two zeroes (extremely rare, 001000000 only)
   E0offset_c0 <= "10000001001"; -- E0 + wE 
   ER_c11 <= E_small_c11(10 downto 0) when small_c11='1'
      else E0offset_c11 - ((10 downto 6 => '0') & E_normal_c11);
   Log_g_c11 <=  Log_small_normd_c11(wF+g-2 downto 0) & "0" when small_c11='1'           -- remove implicit 1
      else Log_normal_normd_c11(targetprec-2 downto targetprec-wF-g-1 );  -- remove implicit 1
   round_c11 <= Log_g_c11(g-1) ; -- sticky is always 1 for a transcendental function 
   -- if round leads to a change of binade, the carry propagation magically updates both mantissa and exponent
   fraX_c11 <= (ER_c11 & Log_g_c11(wF+g-1 downto g)) ; 
   fraY_c11 <= ((wE+wF-1 downto 1 => '0') & round_c11); 
   finalRoundAdder: IntAdder_77_Freq300_uid79
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 Cin => '0',
                 X => fraX_c11,
                 Y => fraY_c11,
                 R => EFR_c11);
   Rexn_c11 <= "110" when ((XExnSgn_c11(2) and (XExnSgn_c11(1) or XExnSgn_c11(0))) or (XExnSgn_c11(1) and XExnSgn_c11(0))) = '1' else
                              "101" when XExnSgn_c11(2 downto 1) = "00"  else
                              "100" when XExnSgn_c11(2 downto 1) = "10"  else
                              "00" & sR_c11 when (((Log_normal_normd_c11(targetprec-1)='0') and (small_c11='0')) or ( (Log_small_normd_c11 (wF+g-1)='0') and (small_c11='1'))) or (ufl_c11 = '1') else
                               "01" & sR_c11;
   R<=  Rexn_c11 & EFR_c11;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid88
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid88 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid88 is
signal Mfull_c12 :  std_logic_vector(40 downto 0);
signal M_c12 :  std_logic_vector(40 downto 0);
signal X_c12 :  std_logic_vector(16 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11, Y_c12 :  std_logic_vector(23 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
            if ce_12 = '1' then
               X_c12 <= X;
               Y_c12 <= Y_c11;
            end if;
         end if;
      end process;
   Mfull_c12 <= std_logic_vector(unsigned(X_c12) * unsigned(Y_c12)); -- multiplier
   M_c12 <= Mfull_c12(40 downto 0);
   R <= M_c12;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid90
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid90 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid90 is
signal Mfull_c12 :  std_logic_vector(40 downto 0);
signal M_c12 :  std_logic_vector(40 downto 0);
signal X_c12 :  std_logic_vector(16 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11, Y_c12 :  std_logic_vector(23 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
            if ce_12 = '1' then
               X_c12 <= X;
               Y_c12 <= Y_c11;
            end if;
         end if;
      end process;
   Mfull_c12 <= std_logic_vector(unsigned(X_c12) * unsigned(Y_c12)); -- multiplier
   M_c12 <= Mfull_c12(40 downto 0);
   R <= M_c12;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x1_Freq300_uid92
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid92 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid92 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x1_Freq300_uid94
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid94 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid94 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (1 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x1_Freq300_uid96
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid96 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid96 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid98
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid98 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid98 is
   component MultTable_Freq300_uid100 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy101_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid100
      port map ( X => Xtable_c11,
                 Y => Y1_copy101_c11);
   Y1_c11 <= Y1_copy101_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid103
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid103 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid103 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid105
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid105 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid105 is
   component MultTable_Freq300_uid107 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy108_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid107
      port map ( X => Xtable_c11,
                 Y => Y1_copy108_c11);
   Y1_c11 <= Y1_copy108_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid110
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid110 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid110 is
   component MultTable_Freq300_uid112 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy113_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid112
      port map ( X => Xtable_c11,
                 Y => Y1_copy113_c11);
   Y1_c11 <= Y1_copy113_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid115
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid115 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid115 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid117
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid117 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid117 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (1 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid119
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid119 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid119 is
   component MultTable_Freq300_uid121 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy122_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid121
      port map ( X => Xtable_c11,
                 Y => Y1_copy122_c11);
   Y1_c11 <= Y1_copy122_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid124
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid124 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid124 is
   component MultTable_Freq300_uid126 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy127_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid126
      port map ( X => Xtable_c11,
                 Y => Y1_copy127_c11);
   Y1_c11 <= Y1_copy127_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid129
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid129 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid129 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid131
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid131 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid131 is
   component MultTable_Freq300_uid133 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy134_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid133
      port map ( X => Xtable_c11,
                 Y => Y1_copy134_c11);
   Y1_c11 <= Y1_copy134_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid136
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid136 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid136 is
   component MultTable_Freq300_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid138
      port map ( X => Xtable_c11,
                 Y => Y1_copy139_c11);
   Y1_c11 <= Y1_copy139_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid141
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid141 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid141 is
   component MultTable_Freq300_uid143 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy144_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid143
      port map ( X => Xtable_c11,
                 Y => Y1_copy144_c11);
   Y1_c11 <= Y1_copy144_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid146
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid146 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid146 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid148
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid148 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid148 is
   component MultTable_Freq300_uid150 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy151_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid150
      port map ( X => Xtable_c11,
                 Y => Y1_copy151_c11);
   Y1_c11 <= Y1_copy151_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid153
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid153 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid153 is
   component MultTable_Freq300_uid155 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy156_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid155
      port map ( X => Xtable_c11,
                 Y => Y1_copy156_c11);
   Y1_c11 <= Y1_copy156_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid158
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid158 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid158 is
   component MultTable_Freq300_uid160 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy161_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid160
      port map ( X => Xtable_c11,
                 Y => Y1_copy161_c11);
   Y1_c11 <= Y1_copy161_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid163
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid163 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid163 is
   component MultTable_Freq300_uid165 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy166_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid165
      port map ( X => Xtable_c11,
                 Y => Y1_copy166_c11);
   Y1_c11 <= Y1_copy166_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid168
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid168 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid168 is
signal Mfull_c12 :  std_logic_vector(40 downto 0);
signal M_c12 :  std_logic_vector(40 downto 0);
signal X_c12 :  std_logic_vector(16 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11, Y_c12 :  std_logic_vector(23 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
            if ce_12 = '1' then
               X_c12 <= X;
               Y_c12 <= Y_c11;
            end if;
         end if;
      end process;
   Mfull_c12 <= std_logic_vector(unsigned(X_c12) * unsigned(Y_c12)); -- multiplier
   M_c12 <= Mfull_c12(40 downto 0);
   R <= M_c12;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid170
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid170 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid170 is
signal Mfull_c12 :  std_logic_vector(40 downto 0);
signal M_c12 :  std_logic_vector(40 downto 0);
signal X_c12 :  std_logic_vector(16 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11, Y_c12 :  std_logic_vector(23 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
            if ce_12 = '1' then
               X_c12 <= X;
               Y_c12 <= Y_c11;
            end if;
         end if;
      end process;
   Mfull_c12 <= std_logic_vector(unsigned(X_c12) * unsigned(Y_c12)); -- multiplier
   M_c12 <= Mfull_c12(40 downto 0);
   R <= M_c12;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid172
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid172 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid172 is
signal Mfull_c12 :  std_logic_vector(40 downto 0);
signal M_c12 :  std_logic_vector(40 downto 0);
signal X_c12 :  std_logic_vector(16 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11, Y_c12 :  std_logic_vector(23 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
            if ce_12 = '1' then
               X_c12 <= X;
               Y_c12 <= Y_c11;
            end if;
         end if;
      end process;
   Mfull_c12 <= std_logic_vector(unsigned(X_c12) * unsigned(Y_c12)); -- multiplier
   M_c12 <= Mfull_c12(40 downto 0);
   R <= M_c12;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid174
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid174 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid174 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid176
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid176 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid176 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid178
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid178 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid178 is
   component MultTable_Freq300_uid180 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy181_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid180
      port map ( X => Xtable_c11,
                 Y => Y1_copy181_c11);
   Y1_c11 <= Y1_copy181_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid183
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid183 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid183 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid185
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid185 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid185 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (1 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid187
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid187 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid187 is
   component MultTable_Freq300_uid189 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy190_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid189
      port map ( X => Xtable_c11,
                 Y => Y1_copy190_c11);
   Y1_c11 <= Y1_copy190_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid192
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid192 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid192 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid194
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid194 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid194 is
   component MultTable_Freq300_uid196 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy197_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid196
      port map ( X => Xtable_c11,
                 Y => Y1_copy197_c11);
   Y1_c11 <= Y1_copy197_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid199
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid199 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid199 is
   component MultTable_Freq300_uid201 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy202_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid201
      port map ( X => Xtable_c11,
                 Y => Y1_copy202_c11);
   Y1_c11 <= Y1_copy202_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid204
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid204 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid204 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid206
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid206 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid206 is
   component MultTable_Freq300_uid208 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy209_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid208
      port map ( X => Xtable_c11,
                 Y => Y1_copy209_c11);
   Y1_c11 <= Y1_copy209_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid211
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid211 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid211 is
   component MultTable_Freq300_uid213 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy214_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid213
      port map ( X => Xtable_c11,
                 Y => Y1_copy214_c11);
   Y1_c11 <= Y1_copy214_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid216
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid216 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid216 is
   component MultTable_Freq300_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid218
      port map ( X => Xtable_c11,
                 Y => Y1_copy219_c11);
   Y1_c11 <= Y1_copy219_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid221
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid221 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid221 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid223
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid223 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid223 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (1 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid225
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid225 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid225 is
   component MultTable_Freq300_uid227 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy228_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid227
      port map ( X => Xtable_c11,
                 Y => Y1_copy228_c11);
   Y1_c11 <= Y1_copy228_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid230
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid230 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid230 is
   component MultTable_Freq300_uid232 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy233_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid232
      port map ( X => Xtable_c11,
                 Y => Y1_copy233_c11);
   Y1_c11 <= Y1_copy233_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid235
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid235 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid235 is
   component MultTable_Freq300_uid237 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy238_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid237
      port map ( X => Xtable_c11,
                 Y => Y1_copy238_c11);
   Y1_c11 <= Y1_copy238_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid240
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid240 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid240 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid242
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid242 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid242 is
   component MultTable_Freq300_uid244 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy245_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid244
      port map ( X => Xtable_c11,
                 Y => Y1_copy245_c11);
   Y1_c11 <= Y1_copy245_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid247
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid247 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid247 is
   component MultTable_Freq300_uid249 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy250_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid249
      port map ( X => Xtable_c11,
                 Y => Y1_copy250_c11);
   Y1_c11 <= Y1_copy250_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid252
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid252 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid252 is
   component MultTable_Freq300_uid254 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy255_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid254
      port map ( X => Xtable_c11,
                 Y => Y1_copy255_c11);
   Y1_c11 <= Y1_copy255_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid257
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid257 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid257 is
   component MultTable_Freq300_uid259 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy260_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid259
      port map ( X => Xtable_c11,
                 Y => Y1_copy260_c11);
   Y1_c11 <= Y1_copy260_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid262
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid262 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid262 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid264
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid264 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid264 is
   component MultTable_Freq300_uid266 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy267_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid266
      port map ( X => Xtable_c11,
                 Y => Y1_copy267_c11);
   Y1_c11 <= Y1_copy267_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid269
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid269 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid269 is
   component MultTable_Freq300_uid271 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy272_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid271
      port map ( X => Xtable_c11,
                 Y => Y1_copy272_c11);
   Y1_c11 <= Y1_copy272_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid274
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid274 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid274 is
   component MultTable_Freq300_uid276 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy277_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid276
      port map ( X => Xtable_c11,
                 Y => Y1_copy277_c11);
   Y1_c11 <= Y1_copy277_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid279
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid279 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid279 is
   component MultTable_Freq300_uid281 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy282_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid281
      port map ( X => Xtable_c11,
                 Y => Y1_copy282_c11);
   Y1_c11 <= Y1_copy282_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid284
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid284 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid284 is
   component MultTable_Freq300_uid286 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy287_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid286
      port map ( X => Xtable_c11,
                 Y => Y1_copy287_c11);
   Y1_c11 <= Y1_copy287_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid289
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid289 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid289 is
signal replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (1 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid291
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid291 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid291 is
   component MultTable_Freq300_uid293 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy294_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid293
      port map ( X => Xtable_c11,
                 Y => Y1_copy294_c11);
   Y1_c11 <= Y1_copy294_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid296
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid296 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid296 is
   component MultTable_Freq300_uid298 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy299_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid298
      port map ( X => Xtable_c11,
                 Y => Y1_copy299_c11);
   Y1_c11 <= Y1_copy299_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid301
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid301 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid301 is
   component MultTable_Freq300_uid303 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy304_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid303
      port map ( X => Xtable_c11,
                 Y => Y1_copy304_c11);
   Y1_c11 <= Y1_copy304_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid306
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid306 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid306 is
   component MultTable_Freq300_uid308 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy309_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid308
      port map ( X => Xtable_c11,
                 Y => Y1_copy309_c11);
   Y1_c11 <= Y1_copy309_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid311
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid311 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid311 is
   component MultTable_Freq300_uid313 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy314_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid313
      port map ( X => Xtable_c11,
                 Y => Y1_copy314_c11);
   Y1_c11 <= Y1_copy314_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid316
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid316 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid316 is
signal replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (1 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid318
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid318 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid318 is
   component MultTable_Freq300_uid320 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy321_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid320
      port map ( X => Xtable_c11,
                 Y => Y1_copy321_c11);
   Y1_c11 <= Y1_copy321_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid323
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid323 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid323 is
   component MultTable_Freq300_uid325 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy326_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid325
      port map ( X => Xtable_c11,
                 Y => Y1_copy326_c11);
   Y1_c11 <= Y1_copy326_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid328
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid328 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid328 is
   component MultTable_Freq300_uid330 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy331_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid330
      port map ( X => Xtable_c11,
                 Y => Y1_copy331_c11);
   Y1_c11 <= Y1_copy331_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid333
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid333 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid333 is
   component MultTable_Freq300_uid335 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy336_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid335
      port map ( X => Xtable_c11,
                 Y => Y1_copy336_c11);
   Y1_c11 <= Y1_copy336_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid338
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid338 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid338 is
   component MultTable_Freq300_uid340 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy341_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid340
      port map ( X => Xtable_c11,
                 Y => Y1_copy341_c11);
   Y1_c11 <= Y1_copy341_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid343
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid343 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid343 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid345
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid345 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid345 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid347
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid347 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid347 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid349
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid349 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid349 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid351
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid351 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid351 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid353
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid353 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid353 is
   component MultTable_Freq300_uid355 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy356_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid355
      port map ( X => Xtable_c11,
                 Y => Y1_copy356_c11);
   Y1_c11 <= Y1_copy356_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid358
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid358 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid358 is
   component MultTable_Freq300_uid360 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy361_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid360
      port map ( X => Xtable_c11,
                 Y => Y1_copy361_c11);
   Y1_c11 <= Y1_copy361_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid363
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid363 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid363 is
   component MultTable_Freq300_uid365 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy366_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid365
      port map ( X => Xtable_c11,
                 Y => Y1_copy366_c11);
   Y1_c11 <= Y1_copy366_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid368
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid368 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid368 is
   component MultTable_Freq300_uid370 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy371_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid370
      port map ( X => Xtable_c11,
                 Y => Y1_copy371_c11);
   Y1_c11 <= Y1_copy371_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid373
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid373 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid373 is
   component MultTable_Freq300_uid375 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy376_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid375
      port map ( X => Xtable_c11,
                 Y => Y1_copy376_c11);
   Y1_c11 <= Y1_copy376_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid378
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid378 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid378 is
   component MultTable_Freq300_uid380 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy381_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid380
      port map ( X => Xtable_c11,
                 Y => Y1_copy381_c11);
   Y1_c11 <= Y1_copy381_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid383
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid383 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid383 is
   component MultTable_Freq300_uid385 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy386_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid385
      port map ( X => Xtable_c11,
                 Y => Y1_copy386_c11);
   Y1_c11 <= Y1_copy386_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid388
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid388 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid388 is
   component MultTable_Freq300_uid390 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy391_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid390
      port map ( X => Xtable_c11,
                 Y => Y1_copy391_c11);
   Y1_c11 <= Y1_copy391_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid393
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid393 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid393 is
   component MultTable_Freq300_uid395 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy396_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid395
      port map ( X => Xtable_c11,
                 Y => Y1_copy396_c11);
   Y1_c11 <= Y1_copy396_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid398
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid398 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid398 is
   component MultTable_Freq300_uid400 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy401_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid400
      port map ( X => Xtable_c11,
                 Y => Y1_copy401_c11);
   Y1_c11 <= Y1_copy401_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid403
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid403 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid403 is
   component MultTable_Freq300_uid405 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy406_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid405
      port map ( X => Xtable_c11,
                 Y => Y1_copy406_c11);
   Y1_c11 <= Y1_copy406_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid408
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid408 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid408 is
   component MultTable_Freq300_uid410 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy411_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid410
      port map ( X => Xtable_c11,
                 Y => Y1_copy411_c11);
   Y1_c11 <= Y1_copy411_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid413
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid413 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid413 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid415
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid415 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid415 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid417
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid417 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid417 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid419
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid419 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid419 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid421
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid421 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid421 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid423
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid423 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid423 is
   component MultTable_Freq300_uid425 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy426_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid425
      port map ( X => Xtable_c11,
                 Y => Y1_copy426_c11);
   Y1_c11 <= Y1_copy426_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid428
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid428 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid428 is
   component MultTable_Freq300_uid430 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy431_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid430
      port map ( X => Xtable_c11,
                 Y => Y1_copy431_c11);
   Y1_c11 <= Y1_copy431_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid433
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid433 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid433 is
   component MultTable_Freq300_uid435 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy436_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid435
      port map ( X => Xtable_c11,
                 Y => Y1_copy436_c11);
   Y1_c11 <= Y1_copy436_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid438
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid438 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid438 is
   component MultTable_Freq300_uid440 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy441_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid440
      port map ( X => Xtable_c11,
                 Y => Y1_copy441_c11);
   Y1_c11 <= Y1_copy441_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid443
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid443 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid443 is
   component MultTable_Freq300_uid445 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy446_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid445
      port map ( X => Xtable_c11,
                 Y => Y1_copy446_c11);
   Y1_c11 <= Y1_copy446_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid448
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid448 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid448 is
   component MultTable_Freq300_uid450 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy451_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid450
      port map ( X => Xtable_c11,
                 Y => Y1_copy451_c11);
   Y1_c11 <= Y1_copy451_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid453
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid453 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid453 is
   component MultTable_Freq300_uid455 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy456_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid455
      port map ( X => Xtable_c11,
                 Y => Y1_copy456_c11);
   Y1_c11 <= Y1_copy456_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid458
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid458 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid458 is
   component MultTable_Freq300_uid460 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy461_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid460
      port map ( X => Xtable_c11,
                 Y => Y1_copy461_c11);
   Y1_c11 <= Y1_copy461_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid463
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid463 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid463 is
   component MultTable_Freq300_uid465 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy466_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid465
      port map ( X => Xtable_c11,
                 Y => Y1_copy466_c11);
   Y1_c11 <= Y1_copy466_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid468
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid468 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid468 is
   component MultTable_Freq300_uid470 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy471_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid470
      port map ( X => Xtable_c11,
                 Y => Y1_copy471_c11);
   Y1_c11 <= Y1_copy471_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid473
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid473 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid473 is
   component MultTable_Freq300_uid475 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy476_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid475
      port map ( X => Xtable_c11,
                 Y => Y1_copy476_c11);
   Y1_c11 <= Y1_copy476_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid478
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid478 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid478 is
   component MultTable_Freq300_uid480 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy481_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid480
      port map ( X => Xtable_c11,
                 Y => Y1_copy481_c11);
   Y1_c11 <= Y1_copy481_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid483
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid483 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid483 is
signal replicated_c11 :  std_logic_vector(0 downto 0);
signal prod_c11 :  std_logic_vector(0 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (0 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid485
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid485 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid485 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid487
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid487 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid487 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid489
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid489 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid489 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid491
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid491 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid491 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid493
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid493 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid493 is
   component MultTable_Freq300_uid495 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy496_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid495
      port map ( X => Xtable_c11,
                 Y => Y1_copy496_c11);
   Y1_c11 <= Y1_copy496_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid498
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid498 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid498 is
   component MultTable_Freq300_uid500 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy501_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid500
      port map ( X => Xtable_c11,
                 Y => Y1_copy501_c11);
   Y1_c11 <= Y1_copy501_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid503
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid503 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid503 is
   component MultTable_Freq300_uid505 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy506_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid505
      port map ( X => Xtable_c11,
                 Y => Y1_copy506_c11);
   Y1_c11 <= Y1_copy506_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid508
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid508 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid508 is
   component MultTable_Freq300_uid510 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy511_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid510
      port map ( X => Xtable_c11,
                 Y => Y1_copy511_c11);
   Y1_c11 <= Y1_copy511_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid513
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid513 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid513 is
   component MultTable_Freq300_uid515 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy516_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid515
      port map ( X => Xtable_c11,
                 Y => Y1_copy516_c11);
   Y1_c11 <= Y1_copy516_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid518
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid518 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid518 is
   component MultTable_Freq300_uid520 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy521_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid520
      port map ( X => Xtable_c11,
                 Y => Y1_copy521_c11);
   Y1_c11 <= Y1_copy521_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid523
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid523 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid523 is
   component MultTable_Freq300_uid525 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(3 downto 0);
signal Y1_c11 :  std_logic_vector(3 downto 0);
signal Y1_copy526_c11 :  std_logic_vector(3 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid525
      port map ( X => Xtable_c11,
                 Y => Y1_copy526_c11);
   Y1_c11 <= Y1_copy526_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid528
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid528 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid528 is
   component MultTable_Freq300_uid530 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy531_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid530
      port map ( X => Xtable_c11,
                 Y => Y1_copy531_c11);
   Y1_c11 <= Y1_copy531_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid533
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid533 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid533 is
   component MultTable_Freq300_uid535 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy536_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid535
      port map ( X => Xtable_c11,
                 Y => Y1_copy536_c11);
   Y1_c11 <= Y1_copy536_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid538
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid538 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid538 is
   component MultTable_Freq300_uid540 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy541_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid540
      port map ( X => Xtable_c11,
                 Y => Y1_copy541_c11);
   Y1_c11 <= Y1_copy541_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid543
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid543 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid543 is
   component MultTable_Freq300_uid545 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy546_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid545
      port map ( X => Xtable_c11,
                 Y => Y1_copy546_c11);
   Y1_c11 <= Y1_copy546_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid548
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid548 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid548 is
   component MultTable_Freq300_uid550 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy551_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid550
      port map ( X => Xtable_c11,
                 Y => Y1_copy551_c11);
   Y1_c11 <= Y1_copy551_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid553
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid553 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid553 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid555
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid555 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid555 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid557
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid557 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid557 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid559
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid559 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid559 is
signal replicated_c0, replicated_c1, replicated_c2, replicated_c3, replicated_c4, replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9, replicated_c10, replicated_c11 :  std_logic_vector(3 downto 0);
signal prod_c11 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               replicated_c1 <= replicated_c0;
            end if;
            if ce_2 = '1' then
               replicated_c2 <= replicated_c1;
            end if;
            if ce_3 = '1' then
               replicated_c3 <= replicated_c2;
            end if;
            if ce_4 = '1' then
               replicated_c4 <= replicated_c3;
            end if;
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
            if ce_10 = '1' then
               replicated_c10 <= replicated_c9;
            end if;
            if ce_11 = '1' then
               replicated_c11 <= replicated_c10;
            end if;
         end if;
      end process;
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c11 <= X and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid561
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid561 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid561 is
signal replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (1 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid563
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid563 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid563 is
   component MultTable_Freq300_uid565 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy566_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid565
      port map ( X => Xtable_c11,
                 Y => Y1_copy566_c11);
   Y1_c11 <= Y1_copy566_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid568
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid568 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid568 is
   component MultTable_Freq300_uid570 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy571_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid570
      port map ( X => Xtable_c11,
                 Y => Y1_copy571_c11);
   Y1_c11 <= Y1_copy571_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid573
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid573 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid573 is
   component MultTable_Freq300_uid575 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy576_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid575
      port map ( X => Xtable_c11,
                 Y => Y1_copy576_c11);
   Y1_c11 <= Y1_copy576_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid578
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid578 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid578 is
   component MultTable_Freq300_uid580 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy581_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid580
      port map ( X => Xtable_c11,
                 Y => Y1_copy581_c11);
   Y1_c11 <= Y1_copy581_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid583
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid583 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid583 is
   component MultTable_Freq300_uid585 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy586_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid585
      port map ( X => Xtable_c11,
                 Y => Y1_copy586_c11);
   Y1_c11 <= Y1_copy586_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid588
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid588 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid588 is
signal replicated_c11 :  std_logic_vector(1 downto 0);
signal prod_c11 :  std_logic_vector(1 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
   replicated_c11 <= (1 downto 0 => X(0));
   prod_c11 <= Y_c11 and replicated_c11;
   R <= prod_c11;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid590
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid590 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid590 is
   component MultTable_Freq300_uid592 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy593_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid592
      port map ( X => Xtable_c11,
                 Y => Y1_copy593_c11);
   Y1_c11 <= Y1_copy593_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid595
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid595 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid595 is
   component MultTable_Freq300_uid597 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy598_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid597
      port map ( X => Xtable_c11,
                 Y => Y1_copy598_c11);
   Y1_c11 <= Y1_copy598_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid600
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid600 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid600 is
   component MultTable_Freq300_uid602 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy603_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid602
      port map ( X => Xtable_c11,
                 Y => Y1_copy603_c11);
   Y1_c11 <= Y1_copy603_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid605
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid605 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid605 is
   component MultTable_Freq300_uid607 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy608_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid607
      port map ( X => Xtable_c11,
                 Y => Y1_copy608_c11);
   Y1_c11 <= Y1_copy608_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid610
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid610 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid610 is
   component MultTable_Freq300_uid612 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c11 :  std_logic_vector(4 downto 0);
signal Y1_c11 :  std_logic_vector(4 downto 0);
signal Y1_copy613_c11 :  std_logic_vector(4 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
            end if;
         end if;
      end process;
Xtable_c11 <= Y_c11 & X;
   R <= Y1_c11;
   TableMult: MultTable_Freq300_uid612
      port map ( X => Xtable_c11,
                 Y => Y1_copy613_c11);
   Y1_c11 <= Y1_copy613_c11; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_75_Freq300_uid1472
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_75_Freq300_uid1472 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
          X : in  std_logic_vector(74 downto 0);
          Y : in  std_logic_vector(74 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(74 downto 0)   );
end entity;

architecture arch of IntAdder_75_Freq300_uid1472 is
signal Rtmp_c14 :  std_logic_vector(74 downto 0);
signal X_c14 :  std_logic_vector(74 downto 0);
signal Y_c14 :  std_logic_vector(74 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               X_c14 <= X;
               Y_c14 <= Y;
               Cin_c14 <= Cin_c13;
            end if;
         end if;
      end process;
   Rtmp_c14 <= X_c14 + Y_c14 + Cin_c14;
   R <= Rtmp_c14;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_67x53_70_Freq300_uid84
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_67x53_70_Freq300_uid84 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
          X : in  std_logic_vector(66 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(69 downto 0)   );
end entity;

architecture arch of IntMultiplier_67x53_70_Freq300_uid84 is
   component DSPBlock_17x24_Freq300_uid88 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid90 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid92 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid94 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid96 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid98 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid103 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid105 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid110 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid115 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid117 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid119 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid124 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid129 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid131 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid136 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid141 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid146 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid148 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid153 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid158 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid163 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid168 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid170 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid172 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid174 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid176 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid178 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid183 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid185 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid187 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid192 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid194 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid199 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid204 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid206 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid211 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid216 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid221 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid223 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid225 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid230 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid235 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid240 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid242 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid247 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid252 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid257 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid262 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid264 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid269 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid274 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid279 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid284 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid289 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid291 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid296 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid301 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid306 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid311 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid316 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid318 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid323 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid328 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid333 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid338 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid343 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid345 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid347 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid349 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid351 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid353 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid358 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid363 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid368 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid373 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid378 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid383 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid388 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid393 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid398 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid403 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid408 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid413 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid415 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid417 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid419 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid421 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid423 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid428 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid433 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid438 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid443 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid448 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid453 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid458 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid463 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid468 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid473 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid478 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid483 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid485 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid487 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid489 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid491 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid493 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid498 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid503 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid508 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid513 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid518 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid523 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid528 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid533 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid538 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid543 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid548 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid553 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid555 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid557 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid559 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid561 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid563 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid568 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid573 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid578 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid583 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid588 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid590 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid595 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid600 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid605 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid610 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid616 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid626 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid650 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid712 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid958 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_75_Freq300_uid1472 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
             X : in  std_logic_vector(74 downto 0);
             Y : in  std_logic_vector(74 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(74 downto 0)   );
   end component;

signal XX_m85_c11 :  std_logic_vector(66 downto 0);
signal YY_m85_c0 :  std_logic_vector(52 downto 0);
signal tile_0_X_c11 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c12 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c12 :  unsigned(40-0 downto 0);
signal bh86_w50_0_c12 :  std_logic;
signal bh86_w51_0_c12 :  std_logic;
signal bh86_w52_0_c12 :  std_logic;
signal bh86_w53_0_c12 :  std_logic;
signal bh86_w54_0_c12 :  std_logic;
signal bh86_w55_0_c12 :  std_logic;
signal bh86_w56_0_c12 :  std_logic;
signal bh86_w57_0_c12 :  std_logic;
signal bh86_w58_0_c12 :  std_logic;
signal bh86_w59_0_c12 :  std_logic;
signal bh86_w60_0_c12 :  std_logic;
signal bh86_w61_0_c12 :  std_logic;
signal bh86_w62_0_c12 :  std_logic;
signal bh86_w63_0_c12 :  std_logic;
signal bh86_w64_0_c12 :  std_logic;
signal bh86_w65_0_c12 :  std_logic;
signal bh86_w66_0_c12 :  std_logic;
signal bh86_w67_0_c12 :  std_logic;
signal bh86_w68_0_c12 :  std_logic;
signal bh86_w69_0_c12 :  std_logic;
signal bh86_w70_0_c12 :  std_logic;
signal bh86_w71_0_c12 :  std_logic;
signal bh86_w72_0_c12 :  std_logic;
signal bh86_w73_0_c12 :  std_logic;
signal bh86_w74_0_c12 :  std_logic;
signal bh86_w75_0_c12 :  std_logic;
signal bh86_w76_0_c12 :  std_logic;
signal bh86_w77_0_c12 :  std_logic;
signal bh86_w78_0_c12 :  std_logic;
signal bh86_w79_0_c12 :  std_logic;
signal bh86_w80_0_c12 :  std_logic;
signal bh86_w81_0_c12 :  std_logic;
signal bh86_w82_0_c12 :  std_logic;
signal bh86_w83_0_c12 :  std_logic;
signal bh86_w84_0_c12 :  std_logic;
signal bh86_w85_0_c12 :  std_logic;
signal bh86_w86_0_c12 :  std_logic;
signal bh86_w87_0_c12 :  std_logic;
signal bh86_w88_0_c12 :  std_logic;
signal bh86_w89_0_c12 :  std_logic;
signal bh86_w90_0_c12 :  std_logic;
signal tile_1_X_c11 :  std_logic_vector(16 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_1_output_c12 :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output_c12 :  unsigned(40-0 downto 0);
signal bh86_w33_0_c12, bh86_w33_0_c13 :  std_logic;
signal bh86_w34_0_c12, bh86_w34_0_c13 :  std_logic;
signal bh86_w35_0_c12, bh86_w35_0_c13 :  std_logic;
signal bh86_w36_0_c12, bh86_w36_0_c13 :  std_logic;
signal bh86_w37_0_c12, bh86_w37_0_c13 :  std_logic;
signal bh86_w38_0_c12, bh86_w38_0_c13 :  std_logic;
signal bh86_w39_0_c12, bh86_w39_0_c13 :  std_logic;
signal bh86_w40_0_c12 :  std_logic;
signal bh86_w41_0_c12 :  std_logic;
signal bh86_w42_0_c12 :  std_logic;
signal bh86_w43_0_c12 :  std_logic;
signal bh86_w44_0_c12 :  std_logic;
signal bh86_w45_0_c12 :  std_logic;
signal bh86_w46_0_c12 :  std_logic;
signal bh86_w47_0_c12 :  std_logic;
signal bh86_w48_0_c12 :  std_logic;
signal bh86_w49_0_c12, bh86_w49_0_c13 :  std_logic;
signal bh86_w50_1_c12, bh86_w50_1_c13 :  std_logic;
signal bh86_w51_1_c12 :  std_logic;
signal bh86_w52_1_c12, bh86_w52_1_c13 :  std_logic;
signal bh86_w53_1_c12 :  std_logic;
signal bh86_w54_1_c12, bh86_w54_1_c13 :  std_logic;
signal bh86_w55_1_c12 :  std_logic;
signal bh86_w56_1_c12 :  std_logic;
signal bh86_w57_1_c12 :  std_logic;
signal bh86_w58_1_c12 :  std_logic;
signal bh86_w59_1_c12 :  std_logic;
signal bh86_w60_1_c12 :  std_logic;
signal bh86_w61_1_c12 :  std_logic;
signal bh86_w62_1_c12 :  std_logic;
signal bh86_w63_1_c12 :  std_logic;
signal bh86_w64_1_c12 :  std_logic;
signal bh86_w65_1_c12 :  std_logic;
signal bh86_w66_1_c12 :  std_logic;
signal bh86_w67_1_c12 :  std_logic;
signal bh86_w68_1_c12 :  std_logic;
signal bh86_w69_1_c12 :  std_logic;
signal bh86_w70_1_c12 :  std_logic;
signal bh86_w71_1_c12 :  std_logic;
signal bh86_w72_1_c12 :  std_logic;
signal bh86_w73_1_c12 :  std_logic;
signal tile_2_X_c11 :  std_logic_vector(0 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_2_output_c11 :  std_logic_vector(0 downto 0);
signal tile_2_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_1_c11 :  std_logic;
signal tile_3_X_c11 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_3_output_c11 :  std_logic_vector(1 downto 0);
signal tile_3_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w44_2_c11 :  std_logic;
signal bh86_w45_1_c11 :  std_logic;
signal tile_4_X_c11 :  std_logic_vector(0 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_4_output_c11 :  std_logic_vector(0 downto 0);
signal tile_4_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_3_c11 :  std_logic;
signal tile_5_X_c11 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_5_output_c11 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w44_4_c11 :  std_logic;
signal bh86_w45_2_c11 :  std_logic;
signal bh86_w46_1_c11 :  std_logic;
signal bh86_w47_1_c11 :  std_logic;
signal bh86_w48_1_c11 :  std_logic;
signal tile_6_X_c11 :  std_logic_vector(0 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_6_output_c11 :  std_logic_vector(0 downto 0);
signal tile_6_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_5_c11 :  std_logic;
signal tile_7_X_c11 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_7_output_c11 :  std_logic_vector(3 downto 0);
signal tile_7_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w44_6_c11 :  std_logic;
signal bh86_w45_3_c11 :  std_logic;
signal bh86_w46_2_c11 :  std_logic;
signal bh86_w47_2_c11 :  std_logic;
signal tile_8_X_c11 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_8_output_c11 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w46_3_c11 :  std_logic;
signal bh86_w47_3_c11 :  std_logic;
signal bh86_w48_2_c11 :  std_logic;
signal bh86_w49_1_c11 :  std_logic;
signal bh86_w50_2_c11 :  std_logic;
signal tile_9_X_c11 :  std_logic_vector(0 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_9_output_c11 :  std_logic_vector(0 downto 0);
signal tile_9_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_7_c11 :  std_logic;
signal tile_10_X_c11 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_10_output_c11 :  std_logic_vector(1 downto 0);
signal tile_10_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w44_8_c11 :  std_logic;
signal bh86_w45_4_c11 :  std_logic;
signal tile_11_X_c11 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_11_output_c11 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w45_5_c11 :  std_logic;
signal bh86_w46_4_c11 :  std_logic;
signal bh86_w47_4_c11 :  std_logic;
signal bh86_w48_3_c11 :  std_logic;
signal bh86_w49_2_c11 :  std_logic;
signal tile_12_X_c11 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_12_output_c11 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w48_4_c11 :  std_logic;
signal bh86_w49_3_c11 :  std_logic;
signal bh86_w50_3_c11 :  std_logic;
signal bh86_w51_2_c11 :  std_logic;
signal bh86_w52_2_c11 :  std_logic;
signal tile_13_X_c11 :  std_logic_vector(0 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_13_output_c11 :  std_logic_vector(0 downto 0);
signal tile_13_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_9_c11 :  std_logic;
signal tile_14_X_c11 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_14_output_c11 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w44_10_c11 :  std_logic;
signal bh86_w45_6_c11 :  std_logic;
signal bh86_w46_5_c11 :  std_logic;
signal bh86_w47_5_c11 :  std_logic;
signal bh86_w48_5_c11 :  std_logic;
signal tile_15_X_c11 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_15_output_c11 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w47_6_c11 :  std_logic;
signal bh86_w48_6_c11 :  std_logic;
signal bh86_w49_4_c11 :  std_logic;
signal bh86_w50_4_c11 :  std_logic;
signal bh86_w51_3_c11 :  std_logic;
signal tile_16_X_c11 :  std_logic_vector(2 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_16_output_c11 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w50_5_c11 :  std_logic;
signal bh86_w51_4_c11 :  std_logic;
signal bh86_w52_3_c11 :  std_logic;
signal bh86_w53_2_c11 :  std_logic;
signal bh86_w54_2_c11 :  std_logic;
signal tile_17_X_c11 :  std_logic_vector(0 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_17_output_c11 :  std_logic_vector(0 downto 0);
signal tile_17_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_11_c11 :  std_logic;
signal tile_18_X_c11 :  std_logic_vector(1 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_18_output_c11 :  std_logic_vector(3 downto 0);
signal tile_18_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w44_12_c11, bh86_w44_12_c12 :  std_logic;
signal bh86_w45_7_c11 :  std_logic;
signal bh86_w46_6_c11 :  std_logic;
signal bh86_w47_7_c11 :  std_logic;
signal tile_19_X_c11 :  std_logic_vector(2 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_19_output_c11 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w46_7_c11, bh86_w46_7_c12 :  std_logic;
signal bh86_w47_8_c11 :  std_logic;
signal bh86_w48_7_c11 :  std_logic;
signal bh86_w49_5_c11 :  std_logic;
signal bh86_w50_6_c11 :  std_logic;
signal tile_20_X_c11 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_20_output_c11 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w49_6_c11 :  std_logic;
signal bh86_w50_7_c11 :  std_logic;
signal bh86_w51_5_c11 :  std_logic;
signal bh86_w52_4_c11 :  std_logic;
signal bh86_w53_3_c11 :  std_logic;
signal tile_21_X_c11 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_21_output_c11 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w52_5_c11 :  std_logic;
signal bh86_w53_4_c11 :  std_logic;
signal bh86_w54_3_c11 :  std_logic;
signal bh86_w55_2_c11 :  std_logic;
signal bh86_w56_2_c11 :  std_logic;
signal tile_22_X_c11 :  std_logic_vector(16 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_22_output_c12 :  std_logic_vector(40 downto 0);
signal tile_22_filtered_output_c12 :  unsigned(40-0 downto 0);
signal bh86_w74_1_c12 :  std_logic;
signal bh86_w75_1_c12 :  std_logic;
signal bh86_w76_1_c12 :  std_logic;
signal bh86_w77_1_c12 :  std_logic;
signal bh86_w78_1_c12 :  std_logic;
signal bh86_w79_1_c12 :  std_logic;
signal bh86_w80_1_c12 :  std_logic;
signal bh86_w81_1_c12 :  std_logic;
signal bh86_w82_1_c12 :  std_logic;
signal bh86_w83_1_c12 :  std_logic;
signal bh86_w84_1_c12 :  std_logic;
signal bh86_w85_1_c12 :  std_logic;
signal bh86_w86_1_c12 :  std_logic;
signal bh86_w87_1_c12 :  std_logic;
signal bh86_w88_1_c12 :  std_logic;
signal bh86_w89_1_c12 :  std_logic;
signal bh86_w90_1_c12 :  std_logic;
signal bh86_w91_0_c12 :  std_logic;
signal bh86_w92_0_c12 :  std_logic;
signal bh86_w93_0_c12 :  std_logic;
signal bh86_w94_0_c12 :  std_logic;
signal bh86_w95_0_c12 :  std_logic;
signal bh86_w96_0_c12 :  std_logic;
signal bh86_w97_0_c12 :  std_logic;
signal bh86_w98_0_c12, bh86_w98_0_c13 :  std_logic;
signal bh86_w99_0_c12 :  std_logic;
signal bh86_w100_0_c12 :  std_logic;
signal bh86_w101_0_c12 :  std_logic;
signal bh86_w102_0_c12 :  std_logic;
signal bh86_w103_0_c12 :  std_logic;
signal bh86_w104_0_c12 :  std_logic;
signal bh86_w105_0_c12 :  std_logic;
signal bh86_w106_0_c12 :  std_logic;
signal bh86_w107_0_c12 :  std_logic;
signal bh86_w108_0_c12 :  std_logic;
signal bh86_w109_0_c12 :  std_logic;
signal bh86_w110_0_c12 :  std_logic;
signal bh86_w111_0_c12 :  std_logic;
signal bh86_w112_0_c12 :  std_logic;
signal bh86_w113_0_c12 :  std_logic;
signal bh86_w114_0_c12 :  std_logic;
signal tile_23_X_c11 :  std_logic_vector(16 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_23_output_c12 :  std_logic_vector(40 downto 0);
signal tile_23_filtered_output_c12 :  unsigned(40-0 downto 0);
signal bh86_w57_2_c12 :  std_logic;
signal bh86_w58_2_c12 :  std_logic;
signal bh86_w59_2_c12 :  std_logic;
signal bh86_w60_2_c12 :  std_logic;
signal bh86_w61_2_c12 :  std_logic;
signal bh86_w62_2_c12 :  std_logic;
signal bh86_w63_2_c12 :  std_logic;
signal bh86_w64_2_c12 :  std_logic;
signal bh86_w65_2_c12 :  std_logic;
signal bh86_w66_2_c12 :  std_logic;
signal bh86_w67_2_c12 :  std_logic;
signal bh86_w68_2_c12 :  std_logic;
signal bh86_w69_2_c12 :  std_logic;
signal bh86_w70_2_c12 :  std_logic;
signal bh86_w71_2_c12 :  std_logic;
signal bh86_w72_2_c12 :  std_logic;
signal bh86_w73_2_c12 :  std_logic;
signal bh86_w74_2_c12 :  std_logic;
signal bh86_w75_2_c12 :  std_logic;
signal bh86_w76_2_c12 :  std_logic;
signal bh86_w77_2_c12 :  std_logic;
signal bh86_w78_2_c12 :  std_logic;
signal bh86_w79_2_c12 :  std_logic;
signal bh86_w80_2_c12 :  std_logic;
signal bh86_w81_2_c12 :  std_logic;
signal bh86_w82_2_c12 :  std_logic;
signal bh86_w83_2_c12 :  std_logic;
signal bh86_w84_2_c12, bh86_w84_2_c13 :  std_logic;
signal bh86_w85_2_c12 :  std_logic;
signal bh86_w86_2_c12, bh86_w86_2_c13 :  std_logic;
signal bh86_w87_2_c12 :  std_logic;
signal bh86_w88_2_c12 :  std_logic;
signal bh86_w89_2_c12 :  std_logic;
signal bh86_w90_2_c12 :  std_logic;
signal bh86_w91_1_c12 :  std_logic;
signal bh86_w92_1_c12 :  std_logic;
signal bh86_w93_1_c12 :  std_logic;
signal bh86_w94_1_c12 :  std_logic;
signal bh86_w95_1_c12 :  std_logic;
signal bh86_w96_1_c12 :  std_logic;
signal bh86_w97_1_c12 :  std_logic;
signal tile_24_X_c11 :  std_logic_vector(16 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_24_output_c12 :  std_logic_vector(40 downto 0);
signal tile_24_filtered_output_c12 :  unsigned(40-0 downto 0);
signal bh86_w40_1_c12 :  std_logic;
signal bh86_w41_1_c12 :  std_logic;
signal bh86_w42_1_c12 :  std_logic;
signal bh86_w43_1_c12 :  std_logic;
signal bh86_w44_13_c12 :  std_logic;
signal bh86_w45_8_c12 :  std_logic;
signal bh86_w46_8_c12 :  std_logic;
signal bh86_w47_9_c12 :  std_logic;
signal bh86_w48_8_c12 :  std_logic;
signal bh86_w49_7_c12 :  std_logic;
signal bh86_w50_8_c12 :  std_logic;
signal bh86_w51_6_c12 :  std_logic;
signal bh86_w52_6_c12 :  std_logic;
signal bh86_w53_5_c12 :  std_logic;
signal bh86_w54_4_c12 :  std_logic;
signal bh86_w55_3_c12 :  std_logic;
signal bh86_w56_3_c12 :  std_logic;
signal bh86_w57_3_c12 :  std_logic;
signal bh86_w58_3_c12 :  std_logic;
signal bh86_w59_3_c12 :  std_logic;
signal bh86_w60_3_c12 :  std_logic;
signal bh86_w61_3_c12 :  std_logic;
signal bh86_w62_3_c12 :  std_logic;
signal bh86_w63_3_c12 :  std_logic;
signal bh86_w64_3_c12 :  std_logic;
signal bh86_w65_3_c12 :  std_logic;
signal bh86_w66_3_c12 :  std_logic;
signal bh86_w67_3_c12 :  std_logic;
signal bh86_w68_3_c12 :  std_logic;
signal bh86_w69_3_c12 :  std_logic;
signal bh86_w70_3_c12 :  std_logic;
signal bh86_w71_3_c12 :  std_logic;
signal bh86_w72_3_c12 :  std_logic;
signal bh86_w73_3_c12 :  std_logic;
signal bh86_w74_3_c12 :  std_logic;
signal bh86_w75_3_c12 :  std_logic;
signal bh86_w76_3_c12 :  std_logic;
signal bh86_w77_3_c12 :  std_logic;
signal bh86_w78_3_c12, bh86_w78_3_c13 :  std_logic;
signal bh86_w79_3_c12, bh86_w79_3_c13 :  std_logic;
signal bh86_w80_3_c12 :  std_logic;
signal tile_25_X_c11 :  std_logic_vector(0 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_25_output_c11 :  std_logic_vector(0 downto 0);
signal tile_25_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_14_c11 :  std_logic;
signal tile_26_X_c11 :  std_logic_vector(0 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_26_output_c11 :  std_logic_vector(0 downto 0);
signal tile_26_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_15_c11 :  std_logic;
signal tile_27_X_c11 :  std_logic_vector(1 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c11 :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w44_16_c11 :  std_logic;
signal bh86_w45_9_c11 :  std_logic;
signal bh86_w46_9_c11 :  std_logic;
signal bh86_w47_10_c11 :  std_logic;
signal tile_28_X_c11 :  std_logic_vector(0 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_28_output_c11 :  std_logic_vector(0 downto 0);
signal tile_28_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_17_c11 :  std_logic;
signal tile_29_X_c11 :  std_logic_vector(1 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_29_output_c11 :  std_logic_vector(1 downto 0);
signal tile_29_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w44_18_c11 :  std_logic;
signal bh86_w45_10_c11 :  std_logic;
signal tile_30_X_c11 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c11 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w45_11_c11 :  std_logic;
signal bh86_w46_10_c11 :  std_logic;
signal bh86_w47_11_c11 :  std_logic;
signal bh86_w48_9_c11 :  std_logic;
signal bh86_w49_8_c11 :  std_logic;
signal tile_31_X_c11 :  std_logic_vector(0 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_31_output_c11 :  std_logic_vector(0 downto 0);
signal tile_31_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_19_c11 :  std_logic;
signal tile_32_X_c11 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c11 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w44_20_c11 :  std_logic;
signal bh86_w45_12_c11 :  std_logic;
signal bh86_w46_11_c11 :  std_logic;
signal bh86_w47_12_c11 :  std_logic;
signal bh86_w48_10_c11 :  std_logic;
signal tile_33_X_c11 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c11 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w47_13_c11 :  std_logic;
signal bh86_w48_11_c11 :  std_logic;
signal bh86_w49_9_c11 :  std_logic;
signal bh86_w50_9_c11 :  std_logic;
signal bh86_w51_7_c11 :  std_logic;
signal tile_34_X_c11 :  std_logic_vector(0 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_34_output_c11 :  std_logic_vector(0 downto 0);
signal tile_34_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_21_c11 :  std_logic;
signal tile_35_X_c11 :  std_logic_vector(1 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c11 :  std_logic_vector(3 downto 0);
signal tile_35_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w44_22_c11 :  std_logic;
signal bh86_w45_13_c11 :  std_logic;
signal bh86_w46_12_c11 :  std_logic;
signal bh86_w47_14_c11 :  std_logic;
signal tile_36_X_c11 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c11 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w46_13_c11 :  std_logic;
signal bh86_w47_15_c11 :  std_logic;
signal bh86_w48_12_c11 :  std_logic;
signal bh86_w49_10_c11 :  std_logic;
signal bh86_w50_10_c11 :  std_logic;
signal tile_37_X_c11 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_37_output_c11 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w49_11_c11 :  std_logic;
signal bh86_w50_11_c11 :  std_logic;
signal bh86_w51_8_c11 :  std_logic;
signal bh86_w52_7_c11 :  std_logic;
signal bh86_w53_6_c11 :  std_logic;
signal tile_38_X_c11 :  std_logic_vector(0 downto 0);
signal tile_38_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_38_output_c11 :  std_logic_vector(0 downto 0);
signal tile_38_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_23_c11 :  std_logic;
signal tile_39_X_c11 :  std_logic_vector(1 downto 0);
signal tile_39_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_39_output_c11 :  std_logic_vector(1 downto 0);
signal tile_39_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w44_24_c11 :  std_logic;
signal bh86_w45_14_c11 :  std_logic;
signal tile_40_X_c11 :  std_logic_vector(2 downto 0);
signal tile_40_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_40_output_c11 :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w45_15_c11 :  std_logic;
signal bh86_w46_14_c11 :  std_logic;
signal bh86_w47_16_c11 :  std_logic;
signal bh86_w48_13_c11 :  std_logic;
signal bh86_w49_12_c11 :  std_logic;
signal tile_41_X_c11 :  std_logic_vector(2 downto 0);
signal tile_41_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_41_output_c11 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w48_14_c11 :  std_logic;
signal bh86_w49_13_c11 :  std_logic;
signal bh86_w50_12_c11 :  std_logic;
signal bh86_w51_9_c11 :  std_logic;
signal bh86_w52_8_c11 :  std_logic;
signal tile_42_X_c11 :  std_logic_vector(2 downto 0);
signal tile_42_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_42_output_c11 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w51_10_c11 :  std_logic;
signal bh86_w52_9_c11 :  std_logic;
signal bh86_w53_7_c11 :  std_logic;
signal bh86_w54_5_c11 :  std_logic;
signal bh86_w55_4_c11 :  std_logic;
signal tile_43_X_c11 :  std_logic_vector(0 downto 0);
signal tile_43_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_43_output_c11 :  std_logic_vector(0 downto 0);
signal tile_43_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_25_c11 :  std_logic;
signal tile_44_X_c11 :  std_logic_vector(2 downto 0);
signal tile_44_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_44_output_c11 :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w44_26_c11 :  std_logic;
signal bh86_w45_16_c11 :  std_logic;
signal bh86_w46_15_c11 :  std_logic;
signal bh86_w47_17_c11 :  std_logic;
signal bh86_w48_15_c11 :  std_logic;
signal tile_45_X_c11 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_45_output_c11 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w47_18_c11 :  std_logic;
signal bh86_w48_16_c11 :  std_logic;
signal bh86_w49_14_c11 :  std_logic;
signal bh86_w50_13_c11 :  std_logic;
signal bh86_w51_11_c11 :  std_logic;
signal tile_46_X_c11 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_46_output_c11 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w50_14_c11 :  std_logic;
signal bh86_w51_12_c11 :  std_logic;
signal bh86_w52_10_c11 :  std_logic;
signal bh86_w53_8_c11 :  std_logic;
signal bh86_w54_6_c11 :  std_logic;
signal tile_47_X_c11 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_47_output_c11 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w53_9_c11 :  std_logic;
signal bh86_w54_7_c11 :  std_logic;
signal bh86_w55_5_c11 :  std_logic;
signal bh86_w56_4_c11 :  std_logic;
signal bh86_w57_4_c11 :  std_logic;
signal tile_48_X_c11 :  std_logic_vector(0 downto 0);
signal tile_48_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_48_output_c11 :  std_logic_vector(0 downto 0);
signal tile_48_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w44_27_c11 :  std_logic;
signal tile_49_X_c11 :  std_logic_vector(1 downto 0);
signal tile_49_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_49_output_c11 :  std_logic_vector(3 downto 0);
signal tile_49_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w44_28_c11 :  std_logic;
signal bh86_w45_17_c11 :  std_logic;
signal bh86_w46_16_c11 :  std_logic;
signal bh86_w47_19_c11 :  std_logic;
signal tile_50_X_c11 :  std_logic_vector(2 downto 0);
signal tile_50_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_50_output_c11 :  std_logic_vector(4 downto 0);
signal tile_50_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w46_17_c11 :  std_logic;
signal bh86_w47_20_c11 :  std_logic;
signal bh86_w48_17_c11 :  std_logic;
signal bh86_w49_15_c11 :  std_logic;
signal bh86_w50_15_c11 :  std_logic;
signal tile_51_X_c11 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_51_output_c11 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w49_16_c11 :  std_logic;
signal bh86_w50_16_c11 :  std_logic;
signal bh86_w51_13_c11 :  std_logic;
signal bh86_w52_11_c11 :  std_logic;
signal bh86_w53_10_c11 :  std_logic;
signal tile_52_X_c11 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_52_output_c11 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w52_12_c11 :  std_logic;
signal bh86_w53_11_c11 :  std_logic;
signal bh86_w54_8_c11 :  std_logic;
signal bh86_w55_6_c11 :  std_logic;
signal bh86_w56_5_c11 :  std_logic;
signal tile_53_X_c11 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_53_output_c11 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w55_7_c11 :  std_logic;
signal bh86_w56_6_c11 :  std_logic;
signal bh86_w57_5_c11 :  std_logic;
signal bh86_w58_4_c11 :  std_logic;
signal bh86_w59_4_c11 :  std_logic;
signal tile_54_X_c11 :  std_logic_vector(0 downto 0);
signal tile_54_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_54_output_c11 :  std_logic_vector(1 downto 0);
signal tile_54_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w44_29_c11 :  std_logic;
signal bh86_w45_18_c11 :  std_logic;
signal tile_55_X_c11 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_55_output_c11 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w45_19_c11 :  std_logic;
signal bh86_w46_18_c11 :  std_logic;
signal bh86_w47_21_c11 :  std_logic;
signal bh86_w48_18_c11 :  std_logic;
signal bh86_w49_17_c11 :  std_logic;
signal tile_56_X_c11 :  std_logic_vector(2 downto 0);
signal tile_56_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_56_output_c11 :  std_logic_vector(4 downto 0);
signal tile_56_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w48_19_c11 :  std_logic;
signal bh86_w49_18_c11 :  std_logic;
signal bh86_w50_17_c11 :  std_logic;
signal bh86_w51_14_c11 :  std_logic;
signal bh86_w52_13_c11, bh86_w52_13_c12 :  std_logic;
signal tile_57_X_c11 :  std_logic_vector(2 downto 0);
signal tile_57_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_57_output_c11 :  std_logic_vector(4 downto 0);
signal tile_57_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w51_15_c11 :  std_logic;
signal bh86_w52_14_c11 :  std_logic;
signal bh86_w53_12_c11 :  std_logic;
signal bh86_w54_9_c11 :  std_logic;
signal bh86_w55_8_c11 :  std_logic;
signal tile_58_X_c11 :  std_logic_vector(2 downto 0);
signal tile_58_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_58_output_c11 :  std_logic_vector(4 downto 0);
signal tile_58_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w54_10_c11 :  std_logic;
signal bh86_w55_9_c11 :  std_logic;
signal bh86_w56_7_c11 :  std_logic;
signal bh86_w57_6_c11 :  std_logic;
signal bh86_w58_5_c11 :  std_logic;
signal tile_59_X_c11 :  std_logic_vector(2 downto 0);
signal tile_59_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_59_output_c11 :  std_logic_vector(4 downto 0);
signal tile_59_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w57_7_c11 :  std_logic;
signal bh86_w58_6_c11 :  std_logic;
signal bh86_w59_5_c11 :  std_logic;
signal bh86_w60_4_c11 :  std_logic;
signal bh86_w61_4_c11 :  std_logic;
signal tile_60_X_c11 :  std_logic_vector(0 downto 0);
signal tile_60_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_60_output_c11 :  std_logic_vector(1 downto 0);
signal tile_60_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w46_19_c11 :  std_logic;
signal bh86_w47_22_c11 :  std_logic;
signal tile_61_X_c11 :  std_logic_vector(2 downto 0);
signal tile_61_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_61_output_c11 :  std_logic_vector(4 downto 0);
signal tile_61_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w47_23_c11 :  std_logic;
signal bh86_w48_20_c11 :  std_logic;
signal bh86_w49_19_c11 :  std_logic;
signal bh86_w50_18_c11 :  std_logic;
signal bh86_w51_16_c11 :  std_logic;
signal tile_62_X_c11 :  std_logic_vector(2 downto 0);
signal tile_62_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_62_output_c11 :  std_logic_vector(4 downto 0);
signal tile_62_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w50_19_c11 :  std_logic;
signal bh86_w51_17_c11 :  std_logic;
signal bh86_w52_15_c11 :  std_logic;
signal bh86_w53_13_c11 :  std_logic;
signal bh86_w54_11_c11 :  std_logic;
signal tile_63_X_c11 :  std_logic_vector(2 downto 0);
signal tile_63_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_63_output_c11 :  std_logic_vector(4 downto 0);
signal tile_63_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w53_14_c11 :  std_logic;
signal bh86_w54_12_c11 :  std_logic;
signal bh86_w55_10_c11 :  std_logic;
signal bh86_w56_8_c11 :  std_logic;
signal bh86_w57_8_c11 :  std_logic;
signal tile_64_X_c11 :  std_logic_vector(2 downto 0);
signal tile_64_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_64_output_c11 :  std_logic_vector(4 downto 0);
signal tile_64_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w56_9_c11 :  std_logic;
signal bh86_w57_9_c11 :  std_logic;
signal bh86_w58_7_c11 :  std_logic;
signal bh86_w59_6_c11 :  std_logic;
signal bh86_w60_5_c11 :  std_logic;
signal tile_65_X_c11 :  std_logic_vector(2 downto 0);
signal tile_65_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_65_output_c11 :  std_logic_vector(4 downto 0);
signal tile_65_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w59_7_c11 :  std_logic;
signal bh86_w60_6_c11 :  std_logic;
signal bh86_w61_5_c11 :  std_logic;
signal bh86_w62_4_c11 :  std_logic;
signal bh86_w63_4_c11 :  std_logic;
signal tile_66_X_c11 :  std_logic_vector(0 downto 0);
signal tile_66_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_66_output_c11 :  std_logic_vector(0 downto 0);
signal tile_66_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w98_1_c11 :  std_logic;
signal tile_67_X_c11 :  std_logic_vector(3 downto 0);
signal tile_67_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_67_output_c11 :  std_logic_vector(3 downto 0);
signal tile_67_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w99_1_c11 :  std_logic;
signal bh86_w100_1_c11 :  std_logic;
signal bh86_w101_1_c11 :  std_logic;
signal bh86_w102_1_c11 :  std_logic;
signal tile_68_X_c11 :  std_logic_vector(3 downto 0);
signal tile_68_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_68_output_c11 :  std_logic_vector(3 downto 0);
signal tile_68_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w103_1_c11 :  std_logic;
signal bh86_w104_1_c11 :  std_logic;
signal bh86_w105_1_c11 :  std_logic;
signal bh86_w106_1_c11 :  std_logic;
signal tile_69_X_c11 :  std_logic_vector(3 downto 0);
signal tile_69_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_69_output_c11 :  std_logic_vector(3 downto 0);
signal tile_69_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w107_1_c11 :  std_logic;
signal bh86_w108_1_c11 :  std_logic;
signal bh86_w109_1_c11 :  std_logic;
signal bh86_w110_1_c11 :  std_logic;
signal tile_70_X_c11 :  std_logic_vector(3 downto 0);
signal tile_70_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_70_output_c11 :  std_logic_vector(3 downto 0);
signal tile_70_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w111_1_c11 :  std_logic;
signal bh86_w112_1_c11 :  std_logic;
signal bh86_w113_1_c11 :  std_logic;
signal bh86_w114_1_c11 :  std_logic;
signal tile_71_X_c11 :  std_logic_vector(1 downto 0);
signal tile_71_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_71_output_c11 :  std_logic_vector(3 downto 0);
signal tile_71_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w99_2_c11 :  std_logic;
signal bh86_w100_2_c11 :  std_logic;
signal bh86_w101_2_c11 :  std_logic;
signal bh86_w102_2_c11 :  std_logic;
signal tile_72_X_c11 :  std_logic_vector(2 downto 0);
signal tile_72_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_72_output_c11 :  std_logic_vector(4 downto 0);
signal tile_72_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w101_3_c11 :  std_logic;
signal bh86_w102_3_c11 :  std_logic;
signal bh86_w103_2_c11 :  std_logic;
signal bh86_w104_2_c11 :  std_logic;
signal bh86_w105_2_c11 :  std_logic;
signal tile_73_X_c11 :  std_logic_vector(2 downto 0);
signal tile_73_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_73_output_c11 :  std_logic_vector(4 downto 0);
signal tile_73_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w104_3_c11 :  std_logic;
signal bh86_w105_3_c11 :  std_logic;
signal bh86_w106_2_c11 :  std_logic;
signal bh86_w107_2_c11 :  std_logic;
signal bh86_w108_2_c11 :  std_logic;
signal tile_74_X_c11 :  std_logic_vector(2 downto 0);
signal tile_74_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_74_output_c11 :  std_logic_vector(4 downto 0);
signal tile_74_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w107_3_c11 :  std_logic;
signal bh86_w108_3_c11 :  std_logic;
signal bh86_w109_2_c11 :  std_logic;
signal bh86_w110_2_c11 :  std_logic;
signal bh86_w111_2_c11 :  std_logic;
signal tile_75_X_c11 :  std_logic_vector(2 downto 0);
signal tile_75_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_75_output_c11 :  std_logic_vector(4 downto 0);
signal tile_75_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w110_3_c11 :  std_logic;
signal bh86_w111_3_c11 :  std_logic;
signal bh86_w112_2_c11 :  std_logic;
signal bh86_w113_2_c11 :  std_logic;
signal bh86_w114_2_c11 :  std_logic;
signal tile_76_X_c11 :  std_logic_vector(2 downto 0);
signal tile_76_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_76_output_c11 :  std_logic_vector(4 downto 0);
signal tile_76_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w113_3_c11 :  std_logic;
signal bh86_w114_3_c11 :  std_logic;
signal bh86_w115_0_c11 :  std_logic;
signal bh86_w116_0_c11 :  std_logic;
signal bh86_w117_0_c11 :  std_logic;
signal tile_77_X_c11 :  std_logic_vector(1 downto 0);
signal tile_77_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_77_output_c11 :  std_logic_vector(3 downto 0);
signal tile_77_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w101_4_c11 :  std_logic;
signal bh86_w102_4_c11 :  std_logic;
signal bh86_w103_3_c11 :  std_logic;
signal bh86_w104_4_c11 :  std_logic;
signal tile_78_X_c11 :  std_logic_vector(2 downto 0);
signal tile_78_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_78_output_c11 :  std_logic_vector(4 downto 0);
signal tile_78_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w103_4_c11 :  std_logic;
signal bh86_w104_5_c11, bh86_w104_5_c12 :  std_logic;
signal bh86_w105_4_c11 :  std_logic;
signal bh86_w106_3_c11 :  std_logic;
signal bh86_w107_4_c11 :  std_logic;
signal tile_79_X_c11 :  std_logic_vector(2 downto 0);
signal tile_79_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_79_output_c11 :  std_logic_vector(4 downto 0);
signal tile_79_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w106_4_c11 :  std_logic;
signal bh86_w107_5_c11 :  std_logic;
signal bh86_w108_4_c11 :  std_logic;
signal bh86_w109_3_c11 :  std_logic;
signal bh86_w110_4_c11 :  std_logic;
signal tile_80_X_c11 :  std_logic_vector(2 downto 0);
signal tile_80_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_80_output_c11 :  std_logic_vector(4 downto 0);
signal tile_80_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w109_4_c11 :  std_logic;
signal bh86_w110_5_c11 :  std_logic;
signal bh86_w111_4_c11 :  std_logic;
signal bh86_w112_3_c11 :  std_logic;
signal bh86_w113_4_c11 :  std_logic;
signal tile_81_X_c11 :  std_logic_vector(2 downto 0);
signal tile_81_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_81_output_c11 :  std_logic_vector(4 downto 0);
signal tile_81_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w112_4_c11 :  std_logic;
signal bh86_w113_5_c11 :  std_logic;
signal bh86_w114_4_c11 :  std_logic;
signal bh86_w115_1_c11 :  std_logic;
signal bh86_w116_1_c11 :  std_logic;
signal tile_82_X_c11 :  std_logic_vector(2 downto 0);
signal tile_82_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_82_output_c11 :  std_logic_vector(4 downto 0);
signal tile_82_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w115_2_c11, bh86_w115_2_c12 :  std_logic;
signal bh86_w116_2_c11 :  std_logic;
signal bh86_w117_1_c11 :  std_logic;
signal bh86_w118_0_c11, bh86_w118_0_c12 :  std_logic;
signal bh86_w119_0_c11 :  std_logic;
signal tile_83_X_c11 :  std_logic_vector(0 downto 0);
signal tile_83_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_83_output_c11 :  std_logic_vector(0 downto 0);
signal tile_83_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w81_3_c11 :  std_logic;
signal tile_84_X_c11 :  std_logic_vector(3 downto 0);
signal tile_84_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_84_output_c11 :  std_logic_vector(3 downto 0);
signal tile_84_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w82_3_c11 :  std_logic;
signal bh86_w83_3_c11 :  std_logic;
signal bh86_w84_3_c11 :  std_logic;
signal bh86_w85_3_c11 :  std_logic;
signal tile_85_X_c11 :  std_logic_vector(3 downto 0);
signal tile_85_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_85_output_c11 :  std_logic_vector(3 downto 0);
signal tile_85_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w86_3_c11 :  std_logic;
signal bh86_w87_3_c11 :  std_logic;
signal bh86_w88_3_c11 :  std_logic;
signal bh86_w89_3_c11 :  std_logic;
signal tile_86_X_c11 :  std_logic_vector(3 downto 0);
signal tile_86_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_86_output_c11 :  std_logic_vector(3 downto 0);
signal tile_86_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w90_3_c11 :  std_logic;
signal bh86_w91_2_c11 :  std_logic;
signal bh86_w92_2_c11 :  std_logic;
signal bh86_w93_2_c11 :  std_logic;
signal tile_87_X_c11 :  std_logic_vector(3 downto 0);
signal tile_87_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_87_output_c11 :  std_logic_vector(3 downto 0);
signal tile_87_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w94_2_c11 :  std_logic;
signal bh86_w95_2_c11 :  std_logic;
signal bh86_w96_2_c11 :  std_logic;
signal bh86_w97_2_c11 :  std_logic;
signal tile_88_X_c11 :  std_logic_vector(1 downto 0);
signal tile_88_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_88_output_c11 :  std_logic_vector(3 downto 0);
signal tile_88_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w82_4_c11 :  std_logic;
signal bh86_w83_4_c11 :  std_logic;
signal bh86_w84_4_c11 :  std_logic;
signal bh86_w85_4_c11 :  std_logic;
signal tile_89_X_c11 :  std_logic_vector(2 downto 0);
signal tile_89_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_89_output_c11 :  std_logic_vector(4 downto 0);
signal tile_89_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w84_5_c11 :  std_logic;
signal bh86_w85_5_c11 :  std_logic;
signal bh86_w86_4_c11 :  std_logic;
signal bh86_w87_4_c11 :  std_logic;
signal bh86_w88_4_c11 :  std_logic;
signal tile_90_X_c11 :  std_logic_vector(2 downto 0);
signal tile_90_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_90_output_c11 :  std_logic_vector(4 downto 0);
signal tile_90_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w87_5_c11 :  std_logic;
signal bh86_w88_5_c11 :  std_logic;
signal bh86_w89_4_c11 :  std_logic;
signal bh86_w90_4_c11 :  std_logic;
signal bh86_w91_3_c11 :  std_logic;
signal tile_91_X_c11 :  std_logic_vector(2 downto 0);
signal tile_91_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_91_output_c11 :  std_logic_vector(4 downto 0);
signal tile_91_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w90_5_c11 :  std_logic;
signal bh86_w91_4_c11 :  std_logic;
signal bh86_w92_3_c11 :  std_logic;
signal bh86_w93_3_c11 :  std_logic;
signal bh86_w94_3_c11 :  std_logic;
signal tile_92_X_c11 :  std_logic_vector(2 downto 0);
signal tile_92_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_92_output_c11 :  std_logic_vector(4 downto 0);
signal tile_92_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w93_4_c11 :  std_logic;
signal bh86_w94_4_c11 :  std_logic;
signal bh86_w95_3_c11 :  std_logic;
signal bh86_w96_3_c11 :  std_logic;
signal bh86_w97_3_c11 :  std_logic;
signal tile_93_X_c11 :  std_logic_vector(2 downto 0);
signal tile_93_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_93_output_c11 :  std_logic_vector(4 downto 0);
signal tile_93_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w96_4_c11 :  std_logic;
signal bh86_w97_4_c11 :  std_logic;
signal bh86_w98_2_c11 :  std_logic;
signal bh86_w99_3_c11 :  std_logic;
signal bh86_w100_3_c11 :  std_logic;
signal tile_94_X_c11 :  std_logic_vector(1 downto 0);
signal tile_94_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_94_output_c11 :  std_logic_vector(3 downto 0);
signal tile_94_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w84_6_c11 :  std_logic;
signal bh86_w85_6_c11 :  std_logic;
signal bh86_w86_5_c11 :  std_logic;
signal bh86_w87_6_c11 :  std_logic;
signal tile_95_X_c11 :  std_logic_vector(2 downto 0);
signal tile_95_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_95_output_c11 :  std_logic_vector(4 downto 0);
signal tile_95_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w86_6_c11 :  std_logic;
signal bh86_w87_7_c11, bh86_w87_7_c12 :  std_logic;
signal bh86_w88_6_c11 :  std_logic;
signal bh86_w89_5_c11 :  std_logic;
signal bh86_w90_6_c11 :  std_logic;
signal tile_96_X_c11 :  std_logic_vector(2 downto 0);
signal tile_96_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_96_output_c11 :  std_logic_vector(4 downto 0);
signal tile_96_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w89_6_c11 :  std_logic;
signal bh86_w90_7_c11 :  std_logic;
signal bh86_w91_5_c11 :  std_logic;
signal bh86_w92_4_c11 :  std_logic;
signal bh86_w93_5_c11 :  std_logic;
signal tile_97_X_c11 :  std_logic_vector(2 downto 0);
signal tile_97_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_97_output_c11 :  std_logic_vector(4 downto 0);
signal tile_97_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w92_5_c11 :  std_logic;
signal bh86_w93_6_c11 :  std_logic;
signal bh86_w94_5_c11 :  std_logic;
signal bh86_w95_4_c11 :  std_logic;
signal bh86_w96_5_c11 :  std_logic;
signal tile_98_X_c11 :  std_logic_vector(2 downto 0);
signal tile_98_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_98_output_c11 :  std_logic_vector(4 downto 0);
signal tile_98_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w95_5_c11 :  std_logic;
signal bh86_w96_6_c11 :  std_logic;
signal bh86_w97_5_c11 :  std_logic;
signal bh86_w98_3_c11 :  std_logic;
signal bh86_w99_4_c11 :  std_logic;
signal tile_99_X_c11 :  std_logic_vector(2 downto 0);
signal tile_99_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_99_output_c11 :  std_logic_vector(4 downto 0);
signal tile_99_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w98_4_c11 :  std_logic;
signal bh86_w99_5_c11 :  std_logic;
signal bh86_w100_4_c11 :  std_logic;
signal bh86_w101_5_c11, bh86_w101_5_c12 :  std_logic;
signal bh86_w102_5_c11 :  std_logic;
signal tile_100_X_c11 :  std_logic_vector(0 downto 0);
signal tile_100_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_100_output_c11 :  std_logic_vector(0 downto 0);
signal tile_100_filtered_output_c11 :  unsigned(0-0 downto 0);
signal bh86_w64_4_c11 :  std_logic;
signal tile_101_X_c11 :  std_logic_vector(3 downto 0);
signal tile_101_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_101_output_c11 :  std_logic_vector(3 downto 0);
signal tile_101_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w65_4_c11 :  std_logic;
signal bh86_w66_4_c11 :  std_logic;
signal bh86_w67_4_c11 :  std_logic;
signal bh86_w68_4_c11 :  std_logic;
signal tile_102_X_c11 :  std_logic_vector(3 downto 0);
signal tile_102_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_102_output_c11 :  std_logic_vector(3 downto 0);
signal tile_102_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w69_4_c11 :  std_logic;
signal bh86_w70_4_c11 :  std_logic;
signal bh86_w71_4_c11 :  std_logic;
signal bh86_w72_4_c11 :  std_logic;
signal tile_103_X_c11 :  std_logic_vector(3 downto 0);
signal tile_103_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_103_output_c11 :  std_logic_vector(3 downto 0);
signal tile_103_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w73_4_c11 :  std_logic;
signal bh86_w74_4_c11 :  std_logic;
signal bh86_w75_4_c11 :  std_logic;
signal bh86_w76_4_c11 :  std_logic;
signal tile_104_X_c11 :  std_logic_vector(3 downto 0);
signal tile_104_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_104_output_c11 :  std_logic_vector(3 downto 0);
signal tile_104_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w77_4_c11 :  std_logic;
signal bh86_w78_4_c11 :  std_logic;
signal bh86_w79_4_c11 :  std_logic;
signal bh86_w80_4_c11 :  std_logic;
signal tile_105_X_c11 :  std_logic_vector(1 downto 0);
signal tile_105_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_105_output_c11 :  std_logic_vector(3 downto 0);
signal tile_105_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w65_5_c11 :  std_logic;
signal bh86_w66_5_c11 :  std_logic;
signal bh86_w67_5_c11 :  std_logic;
signal bh86_w68_5_c11 :  std_logic;
signal tile_106_X_c11 :  std_logic_vector(2 downto 0);
signal tile_106_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_106_output_c11 :  std_logic_vector(4 downto 0);
signal tile_106_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w67_6_c11 :  std_logic;
signal bh86_w68_6_c11 :  std_logic;
signal bh86_w69_5_c11 :  std_logic;
signal bh86_w70_5_c11 :  std_logic;
signal bh86_w71_5_c11 :  std_logic;
signal tile_107_X_c11 :  std_logic_vector(2 downto 0);
signal tile_107_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_107_output_c11 :  std_logic_vector(4 downto 0);
signal tile_107_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w70_6_c11 :  std_logic;
signal bh86_w71_6_c11 :  std_logic;
signal bh86_w72_5_c11 :  std_logic;
signal bh86_w73_5_c11 :  std_logic;
signal bh86_w74_5_c11 :  std_logic;
signal tile_108_X_c11 :  std_logic_vector(2 downto 0);
signal tile_108_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_108_output_c11 :  std_logic_vector(4 downto 0);
signal tile_108_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w73_6_c11 :  std_logic;
signal bh86_w74_6_c11 :  std_logic;
signal bh86_w75_5_c11 :  std_logic;
signal bh86_w76_5_c11 :  std_logic;
signal bh86_w77_5_c11 :  std_logic;
signal tile_109_X_c11 :  std_logic_vector(2 downto 0);
signal tile_109_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_109_output_c11 :  std_logic_vector(4 downto 0);
signal tile_109_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w76_6_c11 :  std_logic;
signal bh86_w77_6_c11 :  std_logic;
signal bh86_w78_5_c11 :  std_logic;
signal bh86_w79_5_c11 :  std_logic;
signal bh86_w80_5_c11 :  std_logic;
signal tile_110_X_c11 :  std_logic_vector(2 downto 0);
signal tile_110_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_110_output_c11 :  std_logic_vector(4 downto 0);
signal tile_110_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w79_6_c11 :  std_logic;
signal bh86_w80_6_c11 :  std_logic;
signal bh86_w81_4_c11 :  std_logic;
signal bh86_w82_5_c11 :  std_logic;
signal bh86_w83_5_c11 :  std_logic;
signal tile_111_X_c11 :  std_logic_vector(1 downto 0);
signal tile_111_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_111_output_c11 :  std_logic_vector(3 downto 0);
signal tile_111_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w67_7_c11 :  std_logic;
signal bh86_w68_7_c11 :  std_logic;
signal bh86_w69_6_c11 :  std_logic;
signal bh86_w70_7_c11 :  std_logic;
signal tile_112_X_c11 :  std_logic_vector(2 downto 0);
signal tile_112_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_112_output_c11 :  std_logic_vector(4 downto 0);
signal tile_112_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w69_7_c11 :  std_logic;
signal bh86_w70_8_c11, bh86_w70_8_c12 :  std_logic;
signal bh86_w71_7_c11 :  std_logic;
signal bh86_w72_6_c11 :  std_logic;
signal bh86_w73_7_c11 :  std_logic;
signal tile_113_X_c11 :  std_logic_vector(2 downto 0);
signal tile_113_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_113_output_c11 :  std_logic_vector(4 downto 0);
signal tile_113_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w72_7_c11 :  std_logic;
signal bh86_w73_8_c11 :  std_logic;
signal bh86_w74_7_c11 :  std_logic;
signal bh86_w75_6_c11 :  std_logic;
signal bh86_w76_7_c11 :  std_logic;
signal tile_114_X_c11 :  std_logic_vector(2 downto 0);
signal tile_114_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_114_output_c11 :  std_logic_vector(4 downto 0);
signal tile_114_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w75_7_c11 :  std_logic;
signal bh86_w76_8_c11 :  std_logic;
signal bh86_w77_7_c11 :  std_logic;
signal bh86_w78_6_c11 :  std_logic;
signal bh86_w79_7_c11 :  std_logic;
signal tile_115_X_c11 :  std_logic_vector(2 downto 0);
signal tile_115_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_115_output_c11 :  std_logic_vector(4 downto 0);
signal tile_115_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w78_7_c11 :  std_logic;
signal bh86_w79_8_c11 :  std_logic;
signal bh86_w80_7_c11 :  std_logic;
signal bh86_w81_5_c11 :  std_logic;
signal bh86_w82_6_c11 :  std_logic;
signal tile_116_X_c11 :  std_logic_vector(2 downto 0);
signal tile_116_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_116_output_c11 :  std_logic_vector(4 downto 0);
signal tile_116_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w81_6_c11 :  std_logic;
signal bh86_w82_7_c11 :  std_logic;
signal bh86_w83_6_c11 :  std_logic;
signal bh86_w84_7_c11, bh86_w84_7_c12 :  std_logic;
signal bh86_w85_7_c11 :  std_logic;
signal tile_117_X_c11 :  std_logic_vector(3 downto 0);
signal tile_117_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_117_output_c11 :  std_logic_vector(3 downto 0);
signal tile_117_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w48_21_c11 :  std_logic;
signal bh86_w49_20_c11 :  std_logic;
signal bh86_w50_20_c11 :  std_logic;
signal bh86_w51_18_c11 :  std_logic;
signal tile_118_X_c11 :  std_logic_vector(3 downto 0);
signal tile_118_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_118_output_c11 :  std_logic_vector(3 downto 0);
signal tile_118_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w52_16_c11 :  std_logic;
signal bh86_w53_15_c11 :  std_logic;
signal bh86_w54_13_c11 :  std_logic;
signal bh86_w55_11_c11 :  std_logic;
signal tile_119_X_c11 :  std_logic_vector(3 downto 0);
signal tile_119_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_119_output_c11 :  std_logic_vector(3 downto 0);
signal tile_119_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w56_10_c11 :  std_logic;
signal bh86_w57_10_c11 :  std_logic;
signal bh86_w58_8_c11 :  std_logic;
signal bh86_w59_8_c11 :  std_logic;
signal tile_120_X_c11 :  std_logic_vector(3 downto 0);
signal tile_120_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_120_output_c11 :  std_logic_vector(3 downto 0);
signal tile_120_filtered_output_c11 :  unsigned(3-0 downto 0);
signal bh86_w60_7_c11 :  std_logic;
signal bh86_w61_6_c11 :  std_logic;
signal bh86_w62_5_c11 :  std_logic;
signal bh86_w63_5_c11 :  std_logic;
signal tile_121_X_c11 :  std_logic_vector(0 downto 0);
signal tile_121_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_121_output_c11 :  std_logic_vector(1 downto 0);
signal tile_121_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w49_21_c11 :  std_logic;
signal bh86_w50_21_c11 :  std_logic;
signal tile_122_X_c11 :  std_logic_vector(2 downto 0);
signal tile_122_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_122_output_c11 :  std_logic_vector(4 downto 0);
signal tile_122_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w50_22_c11 :  std_logic;
signal bh86_w51_19_c11 :  std_logic;
signal bh86_w52_17_c11 :  std_logic;
signal bh86_w53_16_c11 :  std_logic;
signal bh86_w54_14_c11 :  std_logic;
signal tile_123_X_c11 :  std_logic_vector(2 downto 0);
signal tile_123_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_123_output_c11 :  std_logic_vector(4 downto 0);
signal tile_123_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w53_17_c11 :  std_logic;
signal bh86_w54_15_c11 :  std_logic;
signal bh86_w55_12_c11 :  std_logic;
signal bh86_w56_11_c11 :  std_logic;
signal bh86_w57_11_c11 :  std_logic;
signal tile_124_X_c11 :  std_logic_vector(2 downto 0);
signal tile_124_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_124_output_c11 :  std_logic_vector(4 downto 0);
signal tile_124_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w56_12_c11 :  std_logic;
signal bh86_w57_12_c11 :  std_logic;
signal bh86_w58_9_c11 :  std_logic;
signal bh86_w59_9_c11 :  std_logic;
signal bh86_w60_8_c11 :  std_logic;
signal tile_125_X_c11 :  std_logic_vector(2 downto 0);
signal tile_125_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_125_output_c11 :  std_logic_vector(4 downto 0);
signal tile_125_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w59_10_c11 :  std_logic;
signal bh86_w60_9_c11 :  std_logic;
signal bh86_w61_7_c11 :  std_logic;
signal bh86_w62_6_c11 :  std_logic;
signal bh86_w63_6_c11 :  std_logic;
signal tile_126_X_c11 :  std_logic_vector(2 downto 0);
signal tile_126_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_126_output_c11 :  std_logic_vector(4 downto 0);
signal tile_126_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w62_7_c11 :  std_logic;
signal bh86_w63_7_c11 :  std_logic;
signal bh86_w64_5_c11 :  std_logic;
signal bh86_w65_6_c11 :  std_logic;
signal bh86_w66_6_c11 :  std_logic;
signal tile_127_X_c11 :  std_logic_vector(0 downto 0);
signal tile_127_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_127_output_c11 :  std_logic_vector(1 downto 0);
signal tile_127_filtered_output_c11 :  unsigned(1-0 downto 0);
signal bh86_w51_20_c11 :  std_logic;
signal bh86_w52_18_c11 :  std_logic;
signal tile_128_X_c11 :  std_logic_vector(2 downto 0);
signal tile_128_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_128_output_c11 :  std_logic_vector(4 downto 0);
signal tile_128_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w52_19_c11 :  std_logic;
signal bh86_w53_18_c11 :  std_logic;
signal bh86_w54_16_c11 :  std_logic;
signal bh86_w55_13_c11 :  std_logic;
signal bh86_w56_13_c11 :  std_logic;
signal tile_129_X_c11 :  std_logic_vector(2 downto 0);
signal tile_129_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_129_output_c11 :  std_logic_vector(4 downto 0);
signal tile_129_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w55_14_c11 :  std_logic;
signal bh86_w56_14_c11 :  std_logic;
signal bh86_w57_13_c11 :  std_logic;
signal bh86_w58_10_c11 :  std_logic;
signal bh86_w59_11_c11 :  std_logic;
signal tile_130_X_c11 :  std_logic_vector(2 downto 0);
signal tile_130_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_130_output_c11 :  std_logic_vector(4 downto 0);
signal tile_130_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w58_11_c11, bh86_w58_11_c12 :  std_logic;
signal bh86_w59_12_c11 :  std_logic;
signal bh86_w60_10_c11 :  std_logic;
signal bh86_w61_8_c11 :  std_logic;
signal bh86_w62_8_c11 :  std_logic;
signal tile_131_X_c11 :  std_logic_vector(2 downto 0);
signal tile_131_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_131_output_c11 :  std_logic_vector(4 downto 0);
signal tile_131_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w61_9_c11 :  std_logic;
signal bh86_w62_9_c11 :  std_logic;
signal bh86_w63_8_c11, bh86_w63_8_c12 :  std_logic;
signal bh86_w64_6_c11 :  std_logic;
signal bh86_w65_7_c11 :  std_logic;
signal tile_132_X_c11 :  std_logic_vector(2 downto 0);
signal tile_132_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_132_output_c11 :  std_logic_vector(4 downto 0);
signal tile_132_filtered_output_c11 :  unsigned(4-0 downto 0);
signal bh86_w64_7_c11 :  std_logic;
signal bh86_w65_8_c11, bh86_w65_8_c12 :  std_logic;
signal bh86_w66_7_c11 :  std_logic;
signal bh86_w67_8_c11, bh86_w67_8_c12 :  std_logic;
signal bh86_w68_8_c11 :  std_logic;
signal bh86_w44_30_c0, bh86_w44_30_c1, bh86_w44_30_c2, bh86_w44_30_c3, bh86_w44_30_c4, bh86_w44_30_c5, bh86_w44_30_c6, bh86_w44_30_c7, bh86_w44_30_c8, bh86_w44_30_c9, bh86_w44_30_c10, bh86_w44_30_c11 :  std_logic;
signal bh86_w45_20_c0 :  std_logic;
signal bh86_w46_20_c0, bh86_w46_20_c1, bh86_w46_20_c2, bh86_w46_20_c3, bh86_w46_20_c4, bh86_w46_20_c5, bh86_w46_20_c6, bh86_w46_20_c7, bh86_w46_20_c8, bh86_w46_20_c9, bh86_w46_20_c10, bh86_w46_20_c11 :  std_logic;
signal bh86_w47_24_c0, bh86_w47_24_c1, bh86_w47_24_c2, bh86_w47_24_c3, bh86_w47_24_c4, bh86_w47_24_c5, bh86_w47_24_c6, bh86_w47_24_c7, bh86_w47_24_c8, bh86_w47_24_c9, bh86_w47_24_c10, bh86_w47_24_c11 :  std_logic;
signal bh86_w48_22_c0 :  std_logic;
signal bh86_w49_22_c0, bh86_w49_22_c1, bh86_w49_22_c2, bh86_w49_22_c3, bh86_w49_22_c4, bh86_w49_22_c5, bh86_w49_22_c6, bh86_w49_22_c7, bh86_w49_22_c8, bh86_w49_22_c9, bh86_w49_22_c10, bh86_w49_22_c11 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid617_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_31_c12 :  std_logic;
signal bh86_w45_21_c12 :  std_logic;
signal bh86_w46_21_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_copy618_c11, Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_copy618_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid619_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_32_c12 :  std_logic;
signal bh86_w45_22_c12 :  std_logic;
signal bh86_w46_22_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_copy620_c11, Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_copy620_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid621_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_33_c12 :  std_logic;
signal bh86_w45_23_c12 :  std_logic;
signal bh86_w46_23_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_copy622_c11, Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_copy622_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid623_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_34_c12 :  std_logic;
signal bh86_w45_24_c12 :  std_logic;
signal bh86_w46_24_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_copy624_c11, Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_copy624_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid627_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_35_c12 :  std_logic;
signal bh86_w45_25_c12 :  std_logic;
signal bh86_w46_25_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_copy628_c11, Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_copy628_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid629_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w45_26_c12 :  std_logic;
signal bh86_w46_26_c12 :  std_logic;
signal bh86_w47_25_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_copy630_c11, Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_copy630_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid631_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w45_27_c12 :  std_logic;
signal bh86_w46_27_c12 :  std_logic;
signal bh86_w47_26_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_copy632_c11, Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_copy632_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid633_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w45_28_c12 :  std_logic;
signal bh86_w46_28_c12 :  std_logic;
signal bh86_w47_27_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_copy634_c11, Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_copy634_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid635_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_29_c12 :  std_logic;
signal bh86_w47_28_c12 :  std_logic;
signal bh86_w48_23_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_copy636_c11, Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_copy636_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid637_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_30_c12 :  std_logic;
signal bh86_w47_29_c12 :  std_logic;
signal bh86_w48_24_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_copy638_c11, Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_copy638_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid639_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_31_c12 :  std_logic;
signal bh86_w47_30_c12 :  std_logic;
signal bh86_w48_25_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_copy640_c11, Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_copy640_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid641_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_31_c12 :  std_logic;
signal bh86_w48_26_c12 :  std_logic;
signal bh86_w49_23_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_copy642_c11, Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_copy642_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid643_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_32_c12 :  std_logic;
signal bh86_w48_27_c12 :  std_logic;
signal bh86_w49_24_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_copy644_c11, Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_copy644_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid645_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_33_c12 :  std_logic;
signal bh86_w48_28_c12 :  std_logic;
signal bh86_w49_25_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_copy646_c11, Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_copy646_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid647_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_34_c12 :  std_logic;
signal bh86_w48_29_c12 :  std_logic;
signal bh86_w49_26_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_copy648_c11, Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_copy648_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid651_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid651_In1_c11 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_35_c12 :  std_logic;
signal bh86_w48_30_c12 :  std_logic;
signal bh86_w49_27_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_copy652_c11, Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_copy652_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid653_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_31_c12 :  std_logic;
signal bh86_w49_28_c12 :  std_logic;
signal bh86_w50_23_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_copy654_c11, Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_copy654_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid655_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_32_c12 :  std_logic;
signal bh86_w49_29_c12 :  std_logic;
signal bh86_w50_24_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_copy656_c11, Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_copy656_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid657_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_33_c12 :  std_logic;
signal bh86_w49_30_c12 :  std_logic;
signal bh86_w50_25_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_copy658_c11, Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_copy658_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid659_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_31_c12 :  std_logic;
signal bh86_w50_26_c12 :  std_logic;
signal bh86_w51_21_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_copy660_c11, Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_copy660_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid661_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_32_c12 :  std_logic;
signal bh86_w50_27_c12 :  std_logic;
signal bh86_w51_22_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_copy662_c11, Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_copy662_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid663_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_33_c12 :  std_logic;
signal bh86_w50_28_c12 :  std_logic;
signal bh86_w51_23_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_copy664_c11, Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_copy664_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid665_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid665_In1_c11 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_34_c12 :  std_logic;
signal bh86_w50_29_c12 :  std_logic;
signal bh86_w51_24_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_copy666_c11, Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_copy666_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid667_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_30_c12 :  std_logic;
signal bh86_w51_25_c12 :  std_logic;
signal bh86_w52_20_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_copy668_c11, Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_copy668_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid669_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_31_c12 :  std_logic;
signal bh86_w51_26_c12 :  std_logic;
signal bh86_w52_21_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_copy670_c11, Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_copy670_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid671_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_32_c12 :  std_logic;
signal bh86_w51_27_c12 :  std_logic;
signal bh86_w52_22_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_copy672_c11, Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_copy672_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid673_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w51_28_c12 :  std_logic;
signal bh86_w52_23_c12 :  std_logic;
signal bh86_w53_19_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_copy674_c11, Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_copy674_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid675_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w51_29_c12 :  std_logic;
signal bh86_w52_24_c12 :  std_logic;
signal bh86_w53_20_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_copy676_c11, Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_copy676_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid677_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w51_30_c12 :  std_logic;
signal bh86_w52_25_c12 :  std_logic;
signal bh86_w53_21_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_copy678_c11, Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_copy678_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid679_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_26_c12 :  std_logic;
signal bh86_w53_22_c12 :  std_logic;
signal bh86_w54_17_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_copy680_c11, Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_copy680_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid681_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_27_c12 :  std_logic;
signal bh86_w53_23_c12 :  std_logic;
signal bh86_w54_18_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_copy682_c11, Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_copy682_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid683_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid683_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_28_c12 :  std_logic;
signal bh86_w53_24_c12 :  std_logic;
signal bh86_w54_19_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_copy684_c11, Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_copy684_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid685_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_25_c12 :  std_logic;
signal bh86_w54_20_c12 :  std_logic;
signal bh86_w55_15_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_copy686_c11, Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_copy686_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid687_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_26_c12 :  std_logic;
signal bh86_w54_21_c12 :  std_logic;
signal bh86_w55_16_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_copy688_c11, Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_copy688_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid689_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid689_In1_c11 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_27_c12 :  std_logic;
signal bh86_w54_22_c12 :  std_logic;
signal bh86_w55_17_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_copy690_c11, Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_copy690_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid691_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w54_23_c12 :  std_logic;
signal bh86_w55_18_c12 :  std_logic;
signal bh86_w56_15_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_copy692_c11, Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_copy692_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid693_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w54_24_c12 :  std_logic;
signal bh86_w55_19_c12 :  std_logic;
signal bh86_w56_16_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_copy694_c11, Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_copy694_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid695_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w55_20_c12 :  std_logic;
signal bh86_w56_17_c12 :  std_logic;
signal bh86_w57_14_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_copy696_c11, Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_copy696_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid697_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w55_21_c12 :  std_logic;
signal bh86_w56_18_c12 :  std_logic;
signal bh86_w57_15_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_copy698_c11, Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_copy698_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid699_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w56_19_c12 :  std_logic;
signal bh86_w57_16_c12 :  std_logic;
signal bh86_w58_12_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_copy700_c11, Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_copy700_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid701_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w56_20_c12 :  std_logic;
signal bh86_w57_17_c12 :  std_logic;
signal bh86_w58_13_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_copy702_c11, Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_copy702_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid703_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w57_18_c12 :  std_logic;
signal bh86_w58_14_c12 :  std_logic;
signal bh86_w59_13_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_copy704_c11, Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_copy704_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid705_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid705_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w57_19_c12 :  std_logic;
signal bh86_w58_15_c12 :  std_logic;
signal bh86_w59_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_copy706_c11, Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_copy706_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid707_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w58_16_c12 :  std_logic;
signal bh86_w59_15_c12 :  std_logic;
signal bh86_w60_11_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_copy708_c11, Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_copy708_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid709_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w59_16_c12 :  std_logic;
signal bh86_w60_12_c12 :  std_logic;
signal bh86_w61_10_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_copy710_c11, Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_copy710_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid713_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w59_17_c12 :  std_logic;
signal bh86_w60_13_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_copy714_c11, Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_copy714_c12 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid715_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w60_14_c12 :  std_logic;
signal bh86_w61_11_c12 :  std_logic;
signal bh86_w62_10_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_copy716_c11, Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_copy716_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid717_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w61_12_c12 :  std_logic;
signal bh86_w62_11_c12 :  std_logic;
signal bh86_w63_9_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_copy718_c11, Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_copy718_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid719_In0_c11 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w62_12_c12 :  std_logic;
signal bh86_w63_10_c12 :  std_logic;
signal bh86_w64_8_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_copy720_c11, Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_copy720_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid721_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid721_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w63_11_c12 :  std_logic;
signal bh86_w64_9_c12 :  std_logic;
signal bh86_w65_9_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_copy722_c11, Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_copy722_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid723_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w64_10_c12 :  std_logic;
signal bh86_w65_10_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_copy724_c11, Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_copy724_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid725_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid725_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w65_11_c12 :  std_logic;
signal bh86_w66_8_c12 :  std_logic;
signal bh86_w67_9_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_copy726_c11, Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_copy726_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid727_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w66_9_c12 :  std_logic;
signal bh86_w67_10_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_copy728_c11, Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_copy728_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid729_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid729_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w67_11_c12 :  std_logic;
signal bh86_w68_9_c12 :  std_logic;
signal bh86_w69_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_copy730_c11, Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_copy730_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid731_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid731_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w68_10_c12 :  std_logic;
signal bh86_w69_9_c12 :  std_logic;
signal bh86_w70_9_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_copy732_c11, Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_copy732_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid733_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w69_10_c12 :  std_logic;
signal bh86_w70_10_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_copy734_c11, Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_copy734_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid735_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid735_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w70_11_c12 :  std_logic;
signal bh86_w71_8_c12 :  std_logic;
signal bh86_w72_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_copy736_c11, Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_copy736_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid737_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w71_9_c12 :  std_logic;
signal bh86_w72_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_copy738_c11, Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_copy738_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid739_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid739_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w72_10_c12 :  std_logic;
signal bh86_w73_9_c12 :  std_logic;
signal bh86_w74_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_copy740_c11, Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_copy740_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid741_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid741_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w73_10_c12 :  std_logic;
signal bh86_w74_9_c12 :  std_logic;
signal bh86_w75_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_copy742_c11, Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_copy742_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid743_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w74_10_c12 :  std_logic;
signal bh86_w75_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_copy744_c11, Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_copy744_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid745_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid745_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w75_10_c12 :  std_logic;
signal bh86_w76_9_c12 :  std_logic;
signal bh86_w77_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_copy746_c11, Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_copy746_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid747_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid747_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w76_10_c12 :  std_logic;
signal bh86_w77_9_c12 :  std_logic;
signal bh86_w78_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_copy748_c11, Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_copy748_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid749_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w77_10_c12 :  std_logic;
signal bh86_w78_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_copy750_c11, Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_copy750_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid751_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid751_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w78_10_c12 :  std_logic;
signal bh86_w79_9_c12 :  std_logic;
signal bh86_w80_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_copy752_c11, Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_copy752_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid753_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid753_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w79_10_c12 :  std_logic;
signal bh86_w80_9_c12 :  std_logic;
signal bh86_w81_7_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_copy754_c11, Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_copy754_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid755_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w80_10_c12 :  std_logic;
signal bh86_w81_8_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_copy756_c11, Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_copy756_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid757_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid757_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w81_9_c12 :  std_logic;
signal bh86_w82_8_c12 :  std_logic;
signal bh86_w83_7_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_copy758_c11, Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_copy758_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid759_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid759_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w82_9_c12 :  std_logic;
signal bh86_w83_8_c12 :  std_logic;
signal bh86_w84_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_copy760_c11, Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_copy760_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid761_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w83_9_c12 :  std_logic;
signal bh86_w84_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_copy762_c11, Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_copy762_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid763_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid763_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w84_10_c12 :  std_logic;
signal bh86_w85_8_c12 :  std_logic;
signal bh86_w86_7_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_copy764_c11, Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_copy764_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid765_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid765_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w85_9_c12 :  std_logic;
signal bh86_w86_8_c12 :  std_logic;
signal bh86_w87_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_copy766_c11, Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_copy766_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid767_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w86_9_c12 :  std_logic;
signal bh86_w87_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_copy768_c11, Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_copy768_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid769_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid769_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w87_10_c12 :  std_logic;
signal bh86_w88_7_c12 :  std_logic;
signal bh86_w89_7_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_copy770_c11, Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_copy770_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid771_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w88_8_c12 :  std_logic;
signal bh86_w89_8_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_copy772_c11, Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_copy772_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid773_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid773_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w89_9_c12 :  std_logic;
signal bh86_w90_8_c12 :  std_logic;
signal bh86_w91_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_copy774_c11, Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_copy774_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid775_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid775_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w90_9_c12 :  std_logic;
signal bh86_w91_7_c12 :  std_logic;
signal bh86_w92_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_copy776_c11, Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_copy776_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid777_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w91_8_c12 :  std_logic;
signal bh86_w92_7_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_copy778_c11, Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_copy778_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid779_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid779_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w92_8_c12 :  std_logic;
signal bh86_w93_7_c12 :  std_logic;
signal bh86_w94_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_copy780_c11, Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_copy780_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid781_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid781_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w93_8_c12 :  std_logic;
signal bh86_w94_7_c12 :  std_logic;
signal bh86_w95_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_copy782_c11, Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_copy782_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid783_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w94_8_c12 :  std_logic;
signal bh86_w95_7_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_copy784_c11, Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_copy784_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid785_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid785_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w95_8_c12 :  std_logic;
signal bh86_w96_7_c12 :  std_logic;
signal bh86_w97_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_copy786_c11, Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_copy786_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid787_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid787_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w96_8_c12 :  std_logic;
signal bh86_w97_7_c12 :  std_logic;
signal bh86_w98_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_copy788_c11, Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_copy788_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid789_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w97_8_c12 :  std_logic;
signal bh86_w98_6_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_copy790_c11, Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_copy790_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid791_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid791_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w98_7_c12 :  std_logic;
signal bh86_w99_6_c12 :  std_logic;
signal bh86_w100_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_copy792_c11, Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_copy792_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid793_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid793_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w99_7_c12 :  std_logic;
signal bh86_w100_6_c12 :  std_logic;
signal bh86_w101_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_copy794_c11, Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_copy794_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid795_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w100_7_c12 :  std_logic;
signal bh86_w101_7_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_copy796_c11, Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_copy796_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid797_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid797_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w101_8_c12 :  std_logic;
signal bh86_w102_6_c12 :  std_logic;
signal bh86_w103_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_copy798_c11, Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_copy798_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid799_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid799_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w102_7_c12 :  std_logic;
signal bh86_w103_6_c12 :  std_logic;
signal bh86_w104_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_copy800_c11, Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_copy800_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid801_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w103_7_c12 :  std_logic;
signal bh86_w104_7_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_copy802_c11, Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_copy802_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid803_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid803_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w104_8_c12 :  std_logic;
signal bh86_w105_5_c12 :  std_logic;
signal bh86_w106_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_copy804_c11, Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_copy804_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid805_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w105_6_c12 :  std_logic;
signal bh86_w106_6_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_copy806_c11, Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_copy806_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid807_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid807_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w106_7_c12 :  std_logic;
signal bh86_w107_6_c12 :  std_logic;
signal bh86_w108_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_copy808_c11, Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_copy808_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid809_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid809_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w107_7_c12 :  std_logic;
signal bh86_w108_6_c12 :  std_logic;
signal bh86_w109_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_copy810_c11, Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_copy810_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid811_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w108_7_c12 :  std_logic;
signal bh86_w109_6_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_copy812_c11, Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_copy812_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid813_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid813_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w109_7_c12 :  std_logic;
signal bh86_w110_6_c12 :  std_logic;
signal bh86_w111_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_copy814_c11, Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_copy814_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid815_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid815_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w110_7_c12 :  std_logic;
signal bh86_w111_6_c12 :  std_logic;
signal bh86_w112_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_copy816_c11, Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_copy816_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid817_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w111_7_c12 :  std_logic;
signal bh86_w112_6_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_copy818_c11, Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_copy818_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid819_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid819_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w112_7_c12 :  std_logic;
signal bh86_w113_6_c12 :  std_logic;
signal bh86_w114_5_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_copy820_c11, Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_copy820_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid821_In0_c11 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid821_In1_c11 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w113_7_c12 :  std_logic;
signal bh86_w114_6_c12 :  std_logic;
signal bh86_w115_3_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_copy822_c11, Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_copy822_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid823_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid823_In1_c11 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w114_7_c12 :  std_logic;
signal bh86_w115_4_c12 :  std_logic;
signal bh86_w116_3_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_copy824_c11, Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_copy824_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid825_In0_c11 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid825_In1_c11 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w116_4_c12 :  std_logic;
signal bh86_w117_2_c12 :  std_logic;
signal bh86_w118_1_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_copy826_c11, Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_copy826_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid827_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_36_c12 :  std_logic;
signal bh86_w45_29_c12 :  std_logic;
signal bh86_w46_32_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_copy828_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid829_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w45_30_c12 :  std_logic;
signal bh86_w46_33_c12 :  std_logic;
signal bh86_w47_36_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_copy830_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid831_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w45_31_c12 :  std_logic;
signal bh86_w46_34_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_copy832_c12 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid833_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_35_c12 :  std_logic;
signal bh86_w47_37_c12 :  std_logic;
signal bh86_w48_34_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_copy834_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid835_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_36_c12 :  std_logic;
signal bh86_w47_38_c12 :  std_logic;
signal bh86_w48_35_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_copy836_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid837_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_39_c12 :  std_logic;
signal bh86_w48_36_c12 :  std_logic;
signal bh86_w49_35_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_copy838_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid839_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid839_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_40_c12 :  std_logic;
signal bh86_w48_37_c12 :  std_logic;
signal bh86_w49_36_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_copy840_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid841_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_38_c12 :  std_logic;
signal bh86_w49_37_c12 :  std_logic;
signal bh86_w50_33_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_copy842_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid843_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w48_39_c12 :  std_logic;
signal bh86_w49_38_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_copy844_c12 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid845_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_39_c12 :  std_logic;
signal bh86_w50_34_c12 :  std_logic;
signal bh86_w51_31_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_copy846_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid847_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_40_c12 :  std_logic;
signal bh86_w50_35_c12 :  std_logic;
signal bh86_w51_32_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_copy848_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid849_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_36_c12 :  std_logic;
signal bh86_w51_33_c12 :  std_logic;
signal bh86_w52_29_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_copy850_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid851_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid851_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_37_c12 :  std_logic;
signal bh86_w51_34_c12 :  std_logic;
signal bh86_w52_30_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_copy852_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid853_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w51_35_c12 :  std_logic;
signal bh86_w52_31_c12 :  std_logic;
signal bh86_w53_28_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_copy854_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid855_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w51_36_c12 :  std_logic;
signal bh86_w52_32_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_copy856_c12 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid857_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_33_c12 :  std_logic;
signal bh86_w53_29_c12 :  std_logic;
signal bh86_w54_25_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_copy858_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid859_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_34_c12 :  std_logic;
signal bh86_w53_30_c12 :  std_logic;
signal bh86_w54_26_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_copy860_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid861_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_31_c12 :  std_logic;
signal bh86_w54_27_c12 :  std_logic;
signal bh86_w55_22_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_copy862_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid863_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid863_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_32_c12 :  std_logic;
signal bh86_w54_28_c12 :  std_logic;
signal bh86_w55_23_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_copy864_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid865_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w54_29_c12 :  std_logic;
signal bh86_w55_24_c12 :  std_logic;
signal bh86_w56_21_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_copy866_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid867_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w55_25_c12 :  std_logic;
signal bh86_w56_22_c12 :  std_logic;
signal bh86_w57_20_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_copy868_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid869_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w56_23_c12 :  std_logic;
signal bh86_w57_21_c12 :  std_logic;
signal bh86_w58_17_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_copy870_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid871_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w57_22_c12 :  std_logic;
signal bh86_w58_18_c12 :  std_logic;
signal bh86_w59_18_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_copy872_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid873_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w58_19_c12 :  std_logic;
signal bh86_w59_19_c12 :  std_logic;
signal bh86_w60_15_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_copy874_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid875_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid875_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid875_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w59_20_c12 :  std_logic;
signal bh86_w60_16_c12 :  std_logic;
signal bh86_w61_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_copy876_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid877_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w60_17_c12 :  std_logic;
signal bh86_w61_14_c12 :  std_logic;
signal bh86_w62_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_copy878_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid879_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w61_15_c12 :  std_logic;
signal bh86_w62_14_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_copy880_c12 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid881_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w62_15_c12 :  std_logic;
signal bh86_w63_12_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_copy882_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid883_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w63_13_c12 :  std_logic;
signal bh86_w64_11_c12 :  std_logic;
signal bh86_w65_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_copy884_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid885_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w64_12_c12 :  std_logic;
signal bh86_w65_13_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_copy886_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid887_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid887_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w65_14_c12 :  std_logic;
signal bh86_w66_10_c12 :  std_logic;
signal bh86_w67_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_copy888_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid889_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid889_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w67_13_c12 :  std_logic;
signal bh86_w68_11_c12 :  std_logic;
signal bh86_w69_11_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_copy890_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid891_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w69_12_c12 :  std_logic;
signal bh86_w70_12_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_copy892_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid893_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid893_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w70_13_c12 :  std_logic;
signal bh86_w71_10_c12 :  std_logic;
signal bh86_w72_11_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_copy894_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid895_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid895_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w72_12_c12 :  std_logic;
signal bh86_w73_11_c12 :  std_logic;
signal bh86_w74_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_copy896_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid897_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w74_12_c12 :  std_logic;
signal bh86_w75_11_c12 :  std_logic;
signal bh86_w76_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_copy898_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid899_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid899_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w75_12_c12 :  std_logic;
signal bh86_w76_12_c12 :  std_logic;
signal bh86_w77_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_copy900_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid901_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w77_12_c12 :  std_logic;
signal bh86_w78_11_c12 :  std_logic;
signal bh86_w79_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_copy902_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid903_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid903_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w78_12_c12 :  std_logic;
signal bh86_w79_12_c12 :  std_logic;
signal bh86_w80_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_copy904_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid905_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w80_12_c12 :  std_logic;
signal bh86_w81_10_c12 :  std_logic;
signal bh86_w82_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_copy906_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid907_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid907_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w81_11_c12 :  std_logic;
signal bh86_w82_11_c12 :  std_logic;
signal bh86_w83_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_copy908_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid909_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w83_11_c12 :  std_logic;
signal bh86_w84_11_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_copy910_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid911_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid911_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w84_12_c12 :  std_logic;
signal bh86_w85_10_c12 :  std_logic;
signal bh86_w86_10_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_copy912_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid913_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w86_11_c12 :  std_logic;
signal bh86_w87_11_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_copy914_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid915_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid915_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w87_12_c12 :  std_logic;
signal bh86_w88_9_c12 :  std_logic;
signal bh86_w89_10_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_copy916_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid917_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid917_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w89_11_c12 :  std_logic;
signal bh86_w90_10_c12 :  std_logic;
signal bh86_w91_9_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_copy918_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid919_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w91_10_c12 :  std_logic;
signal bh86_w92_9_c12 :  std_logic;
signal bh86_w93_9_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_copy920_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid921_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid921_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w92_10_c12 :  std_logic;
signal bh86_w93_10_c12 :  std_logic;
signal bh86_w94_9_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_copy922_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid923_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w94_10_c12 :  std_logic;
signal bh86_w95_9_c12 :  std_logic;
signal bh86_w96_9_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_copy924_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid925_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid925_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w95_10_c12 :  std_logic;
signal bh86_w96_10_c12 :  std_logic;
signal bh86_w97_9_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_copy926_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid927_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w97_10_c12 :  std_logic;
signal bh86_w98_8_c12 :  std_logic;
signal bh86_w99_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_copy928_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid929_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid929_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w98_9_c12 :  std_logic;
signal bh86_w99_9_c12 :  std_logic;
signal bh86_w100_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_copy930_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid931_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w100_9_c12 :  std_logic;
signal bh86_w101_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_copy932_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid933_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid933_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w101_10_c12 :  std_logic;
signal bh86_w102_8_c12 :  std_logic;
signal bh86_w103_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_copy934_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid935_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w103_9_c12 :  std_logic;
signal bh86_w104_9_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_copy936_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid937_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid937_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w104_10_c12 :  std_logic;
signal bh86_w105_7_c12 :  std_logic;
signal bh86_w106_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_copy938_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid939_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid939_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w106_9_c12 :  std_logic;
signal bh86_w107_8_c12 :  std_logic;
signal bh86_w108_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_copy940_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid941_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w108_9_c12 :  std_logic;
signal bh86_w109_8_c12 :  std_logic;
signal bh86_w110_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_copy942_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid943_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid943_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w109_9_c12 :  std_logic;
signal bh86_w110_9_c12 :  std_logic;
signal bh86_w111_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_copy944_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid945_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w111_9_c12 :  std_logic;
signal bh86_w112_8_c12 :  std_logic;
signal bh86_w113_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_copy946_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid947_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid947_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w112_9_c12 :  std_logic;
signal bh86_w113_9_c12 :  std_logic;
signal bh86_w114_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_copy948_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid949_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid949_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w114_9_c12 :  std_logic;
signal bh86_w115_5_c12 :  std_logic;
signal bh86_w116_5_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_copy950_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid951_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid951_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w116_6_c12 :  std_logic;
signal bh86_w117_3_c12 :  std_logic;
signal bh86_w118_2_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_copy952_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid953_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid953_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid953_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w118_3_c12 :  std_logic;
signal bh86_w119_1_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_copy954_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid955_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w45_32_c12 :  std_logic;
signal bh86_w46_37_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_copy956_c12 :  std_logic_vector(1 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid959_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_38_c12 :  std_logic;
signal bh86_w47_41_c12 :  std_logic;
signal bh86_w48_40_c12 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_copy960_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid961_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w47_42_c12 :  std_logic;
signal bh86_w48_41_c12 :  std_logic;
signal bh86_w49_41_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_copy962_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid963_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_42_c12 :  std_logic;
signal bh86_w49_42_c12 :  std_logic;
signal bh86_w50_38_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_copy964_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid965_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w49_43_c12 :  std_logic;
signal bh86_w50_39_c12 :  std_logic;
signal bh86_w51_37_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_copy966_c12 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid967_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_40_c12 :  std_logic;
signal bh86_w51_38_c12 :  std_logic;
signal bh86_w52_35_c12 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_copy968_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid969_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w51_39_c12 :  std_logic;
signal bh86_w52_36_c12 :  std_logic;
signal bh86_w53_33_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_copy970_c12 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid971_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_37_c12 :  std_logic;
signal bh86_w53_34_c12 :  std_logic;
signal bh86_w54_30_c12 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_copy972_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid973_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid973_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_35_c12 :  std_logic;
signal bh86_w54_31_c12 :  std_logic;
signal bh86_w55_26_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_copy974_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid975_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid975_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w54_32_c12 :  std_logic;
signal bh86_w55_27_c12 :  std_logic;
signal bh86_w56_24_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_copy976_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid977_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w55_28_c12 :  std_logic;
signal bh86_w56_25_c12 :  std_logic;
signal bh86_w57_23_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_copy978_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid979_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w56_26_c12 :  std_logic;
signal bh86_w57_24_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_copy980_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid981_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid981_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w57_25_c12 :  std_logic;
signal bh86_w58_20_c12 :  std_logic;
signal bh86_w59_21_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_copy982_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid983_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w59_22_c12 :  std_logic;
signal bh86_w60_18_c12 :  std_logic;
signal bh86_w61_16_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_copy984_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid985_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w60_19_c12 :  std_logic;
signal bh86_w61_17_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_copy986_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid987_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid987_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w61_18_c12 :  std_logic;
signal bh86_w62_16_c12 :  std_logic;
signal bh86_w63_14_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_copy988_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid989_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid989_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w63_15_c12 :  std_logic;
signal bh86_w64_13_c12 :  std_logic;
signal bh86_w65_15_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_copy990_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid991_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid991_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w65_16_c12 :  std_logic;
signal bh86_w66_11_c12 :  std_logic;
signal bh86_w67_14_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_copy992_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid993_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid993_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w67_15_c12 :  std_logic;
signal bh86_w68_12_c12 :  std_logic;
signal bh86_w69_13_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_copy994_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid995_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid995_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w69_14_c12 :  std_logic;
signal bh86_w70_14_c12 :  std_logic;
signal bh86_w71_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_copy996_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid997_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid997_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w71_12_c12 :  std_logic;
signal bh86_w72_13_c12 :  std_logic;
signal bh86_w73_12_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_copy998_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid999_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid999_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w74_13_c12 :  std_logic;
signal bh86_w75_13_c12 :  std_logic;
signal bh86_w76_13_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_copy1000_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1001_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1001_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w76_14_c12 :  std_logic;
signal bh86_w77_13_c12 :  std_logic;
signal bh86_w78_13_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_copy1002_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1003_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1003_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w78_14_c12 :  std_logic;
signal bh86_w79_13_c12 :  std_logic;
signal bh86_w80_13_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_copy1004_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1005_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1005_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w80_14_c12 :  std_logic;
signal bh86_w81_12_c12 :  std_logic;
signal bh86_w82_12_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_copy1006_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1007_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1007_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w82_13_c12 :  std_logic;
signal bh86_w83_12_c12 :  std_logic;
signal bh86_w84_13_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_copy1008_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1009_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1009_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w84_14_c12 :  std_logic;
signal bh86_w85_11_c12 :  std_logic;
signal bh86_w86_12_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_copy1010_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1011_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1011_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w86_13_c12 :  std_logic;
signal bh86_w87_13_c12 :  std_logic;
signal bh86_w88_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_copy1012_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1013_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1013_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w88_11_c12 :  std_logic;
signal bh86_w89_12_c12 :  std_logic;
signal bh86_w90_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_copy1014_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1015_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1015_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w91_11_c12 :  std_logic;
signal bh86_w92_11_c12 :  std_logic;
signal bh86_w93_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_copy1016_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1017_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1017_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w93_12_c12 :  std_logic;
signal bh86_w94_11_c12 :  std_logic;
signal bh86_w95_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_copy1018_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1019_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1019_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w95_12_c12 :  std_logic;
signal bh86_w96_11_c12 :  std_logic;
signal bh86_w97_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_copy1020_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1021_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1021_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w97_12_c12 :  std_logic;
signal bh86_w98_10_c12 :  std_logic;
signal bh86_w99_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_copy1022_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1023_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1023_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w99_11_c12 :  std_logic;
signal bh86_w100_10_c12 :  std_logic;
signal bh86_w101_11_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_copy1024_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1025_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1025_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w101_12_c12 :  std_logic;
signal bh86_w102_9_c12 :  std_logic;
signal bh86_w103_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_copy1026_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1027_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1027_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w103_11_c12 :  std_logic;
signal bh86_w104_11_c12 :  std_logic;
signal bh86_w105_8_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_copy1028_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1029_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1029_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w105_9_c12 :  std_logic;
signal bh86_w106_10_c12 :  std_logic;
signal bh86_w107_9_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_copy1030_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1031_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1031_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w108_10_c12 :  std_logic;
signal bh86_w109_10_c12 :  std_logic;
signal bh86_w110_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_copy1032_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1033_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1033_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w110_11_c12 :  std_logic;
signal bh86_w111_10_c12 :  std_logic;
signal bh86_w112_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_copy1034_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1035_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1035_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w112_11_c12 :  std_logic;
signal bh86_w113_10_c12 :  std_logic;
signal bh86_w114_10_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_copy1036_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1037_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1037_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w114_11_c12 :  std_logic;
signal bh86_w115_6_c12 :  std_logic;
signal bh86_w116_7_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_copy1038_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1039_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1039_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w116_8_c12 :  std_logic;
signal bh86_w117_4_c12 :  std_logic;
signal bh86_w118_4_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_copy1040_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1041_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1041_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w118_5_c12 :  std_logic;
signal bh86_w119_2_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_copy1042_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1043_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1043_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_39_c12 :  std_logic;
signal bh86_w47_43_c12 :  std_logic;
signal bh86_w48_43_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_copy1044_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1045_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_44_c12 :  std_logic;
signal bh86_w49_44_c12 :  std_logic;
signal bh86_w50_41_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_copy1046_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1047_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w49_45_c12 :  std_logic;
signal bh86_w50_42_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_copy1048_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1049_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1049_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_43_c12 :  std_logic;
signal bh86_w51_40_c12 :  std_logic;
signal bh86_w52_38_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_copy1050_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1051_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w52_39_c12 :  std_logic;
signal bh86_w53_36_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_copy1052_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1053_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w53_37_c12 :  std_logic;
signal bh86_w54_33_c12 :  std_logic;
signal bh86_w55_29_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_copy1054_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1055_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w54_34_c12 :  std_logic;
signal bh86_w55_30_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_copy1056_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1057_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1057_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w55_31_c12 :  std_logic;
signal bh86_w56_27_c12 :  std_logic;
signal bh86_w57_26_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_copy1058_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1059_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1059_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w57_27_c12 :  std_logic;
signal bh86_w58_21_c12 :  std_logic;
signal bh86_w59_23_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_copy1060_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1061_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1061_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w59_24_c12 :  std_logic;
signal bh86_w60_20_c12 :  std_logic;
signal bh86_w61_19_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_copy1062_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1063_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1063_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w61_20_c12 :  std_logic;
signal bh86_w62_17_c12 :  std_logic;
signal bh86_w63_16_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_copy1064_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1065_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1065_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w63_17_c12 :  std_logic;
signal bh86_w64_14_c12 :  std_logic;
signal bh86_w65_17_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_copy1066_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1067_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1067_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w65_18_c12 :  std_logic;
signal bh86_w66_12_c12 :  std_logic;
signal bh86_w67_16_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_copy1068_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1069_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1069_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w67_17_c12 :  std_logic;
signal bh86_w68_13_c12 :  std_logic;
signal bh86_w69_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_copy1070_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1071_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1071_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w69_16_c12 :  std_logic;
signal bh86_w70_15_c12 :  std_logic;
signal bh86_w71_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_copy1072_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1073_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1073_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w71_14_c12 :  std_logic;
signal bh86_w72_14_c12 :  std_logic;
signal bh86_w73_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_copy1074_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1075_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1075_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w73_14_c12 :  std_logic;
signal bh86_w74_14_c12 :  std_logic;
signal bh86_w75_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_copy1076_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1077_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1077_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w76_15_c12 :  std_logic;
signal bh86_w77_14_c12 :  std_logic;
signal bh86_w78_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_copy1078_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1079_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1079_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w78_16_c12 :  std_logic;
signal bh86_w79_14_c12 :  std_logic;
signal bh86_w80_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_copy1080_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1081_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1081_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w80_16_c12 :  std_logic;
signal bh86_w81_13_c12 :  std_logic;
signal bh86_w82_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_copy1082_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1083_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1083_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w82_15_c12 :  std_logic;
signal bh86_w83_13_c12 :  std_logic;
signal bh86_w84_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_copy1084_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1085_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1085_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w84_16_c12 :  std_logic;
signal bh86_w85_12_c12 :  std_logic;
signal bh86_w86_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_copy1086_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1087_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1087_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w86_15_c12 :  std_logic;
signal bh86_w87_14_c12 :  std_logic;
signal bh86_w88_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_copy1088_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1089_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1089_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w88_13_c12 :  std_logic;
signal bh86_w89_13_c12 :  std_logic;
signal bh86_w90_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_copy1090_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1091_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1091_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w90_13_c12 :  std_logic;
signal bh86_w91_12_c12 :  std_logic;
signal bh86_w92_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_copy1092_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1093_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1093_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w93_13_c12 :  std_logic;
signal bh86_w94_12_c12 :  std_logic;
signal bh86_w95_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_copy1094_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1095_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1095_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w95_14_c12 :  std_logic;
signal bh86_w96_12_c12 :  std_logic;
signal bh86_w97_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_copy1096_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1097_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1097_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w97_14_c12 :  std_logic;
signal bh86_w98_11_c12 :  std_logic;
signal bh86_w99_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_copy1098_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1099_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1099_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w99_13_c12 :  std_logic;
signal bh86_w100_11_c12 :  std_logic;
signal bh86_w101_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_copy1100_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1101_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1101_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w101_14_c12 :  std_logic;
signal bh86_w102_10_c12 :  std_logic;
signal bh86_w103_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_copy1102_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1103_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1103_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w103_13_c12 :  std_logic;
signal bh86_w104_12_c12 :  std_logic;
signal bh86_w105_10_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_copy1104_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1105_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1105_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w105_11_c12 :  std_logic;
signal bh86_w106_11_c12 :  std_logic;
signal bh86_w107_10_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_copy1106_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1107_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1107_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w107_11_c12 :  std_logic;
signal bh86_w108_11_c12 :  std_logic;
signal bh86_w109_11_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_copy1108_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1109_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1109_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w110_12_c12 :  std_logic;
signal bh86_w111_11_c12 :  std_logic;
signal bh86_w112_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_copy1110_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1111_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1111_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w112_13_c12 :  std_logic;
signal bh86_w113_11_c12 :  std_logic;
signal bh86_w114_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_copy1112_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1113_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1113_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w114_13_c12 :  std_logic;
signal bh86_w115_7_c12 :  std_logic;
signal bh86_w116_9_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_copy1114_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1115_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1115_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w116_10_c12 :  std_logic;
signal bh86_w117_5_c12 :  std_logic;
signal bh86_w118_6_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_copy1116_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1117_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1117_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w118_7_c12 :  std_logic;
signal bh86_w119_3_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_copy1118_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1119_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1119_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w48_45_c12 :  std_logic;
signal bh86_w49_46_c12 :  std_logic;
signal bh86_w50_44_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_copy1120_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1121_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1121_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w50_45_c12 :  std_logic;
signal bh86_w51_41_c12 :  std_logic;
signal bh86_w52_40_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_copy1122_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1123_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1123_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w52_41_c12 :  std_logic;
signal bh86_w53_38_c12 :  std_logic;
signal bh86_w54_35_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_copy1124_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1125_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w54_36_c12 :  std_logic;
signal bh86_w55_32_c12 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_copy1126_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1127_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1127_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w55_33_c12 :  std_logic;
signal bh86_w56_28_c12 :  std_logic;
signal bh86_w57_28_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_copy1128_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1129_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1129_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w57_29_c12 :  std_logic;
signal bh86_w58_22_c12 :  std_logic;
signal bh86_w59_25_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_copy1130_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1131_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1131_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w59_26_c12 :  std_logic;
signal bh86_w60_21_c12 :  std_logic;
signal bh86_w61_21_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_copy1132_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1133_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1133_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w61_22_c12 :  std_logic;
signal bh86_w62_18_c12 :  std_logic;
signal bh86_w63_18_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_copy1134_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1135_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1135_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w63_19_c12 :  std_logic;
signal bh86_w64_15_c12 :  std_logic;
signal bh86_w65_19_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_copy1136_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1137_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1137_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w65_20_c12 :  std_logic;
signal bh86_w66_13_c12 :  std_logic;
signal bh86_w67_18_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_copy1138_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1139_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1139_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w67_19_c12 :  std_logic;
signal bh86_w68_14_c12 :  std_logic;
signal bh86_w69_17_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_copy1140_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1141_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1141_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w69_18_c12 :  std_logic;
signal bh86_w70_16_c12 :  std_logic;
signal bh86_w71_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_copy1142_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1143_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1143_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w71_16_c12 :  std_logic;
signal bh86_w72_15_c12 :  std_logic;
signal bh86_w73_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_copy1144_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1145_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1145_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w73_16_c12 :  std_logic;
signal bh86_w74_15_c12 :  std_logic;
signal bh86_w75_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_copy1146_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1147_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1147_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w75_16_c12 :  std_logic;
signal bh86_w76_16_c12 :  std_logic;
signal bh86_w77_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_copy1148_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1149_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1149_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w78_17_c12 :  std_logic;
signal bh86_w79_15_c12 :  std_logic;
signal bh86_w80_17_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_copy1150_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1151_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1151_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w80_18_c12 :  std_logic;
signal bh86_w81_14_c12 :  std_logic;
signal bh86_w82_16_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_copy1152_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1153_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1153_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w82_17_c12 :  std_logic;
signal bh86_w83_14_c12 :  std_logic;
signal bh86_w84_17_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_copy1154_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1155_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1155_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w84_18_c12 :  std_logic;
signal bh86_w85_13_c12 :  std_logic;
signal bh86_w86_16_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_copy1156_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1157_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1157_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w86_17_c12 :  std_logic;
signal bh86_w87_15_c12 :  std_logic;
signal bh86_w88_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_copy1158_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1159_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1159_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w88_15_c12, bh86_w88_15_c13 :  std_logic;
signal bh86_w89_14_c12 :  std_logic;
signal bh86_w90_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_copy1160_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1161_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1161_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w90_15_c12 :  std_logic;
signal bh86_w91_13_c12 :  std_logic;
signal bh86_w92_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_copy1162_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1163_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1163_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w92_14_c12 :  std_logic;
signal bh86_w93_14_c12 :  std_logic;
signal bh86_w94_13_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_copy1164_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1165_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1165_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w95_15_c12 :  std_logic;
signal bh86_w96_13_c12 :  std_logic;
signal bh86_w97_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_copy1166_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1167_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1167_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w97_16_c12 :  std_logic;
signal bh86_w98_12_c12 :  std_logic;
signal bh86_w99_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_copy1168_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1169_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1169_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w99_15_c12 :  std_logic;
signal bh86_w100_12_c12 :  std_logic;
signal bh86_w101_15_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_copy1170_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1171_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1171_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w101_16_c12 :  std_logic;
signal bh86_w102_11_c12 :  std_logic;
signal bh86_w103_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_copy1172_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1173_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1173_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w103_15_c12 :  std_logic;
signal bh86_w104_13_c12 :  std_logic;
signal bh86_w105_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_copy1174_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1175_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1175_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w105_13_c12 :  std_logic;
signal bh86_w106_12_c12 :  std_logic;
signal bh86_w107_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_copy1176_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1177_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1177_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w107_13_c12 :  std_logic;
signal bh86_w108_12_c12 :  std_logic;
signal bh86_w109_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_copy1178_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1179_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1179_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w109_13_c12 :  std_logic;
signal bh86_w110_13_c12 :  std_logic;
signal bh86_w111_12_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_copy1180_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1181_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1181_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w112_14_c12 :  std_logic;
signal bh86_w113_12_c12 :  std_logic;
signal bh86_w114_14_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_copy1182_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1183_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1183_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w114_15_c12 :  std_logic;
signal bh86_w115_8_c12, bh86_w115_8_c13 :  std_logic;
signal bh86_w116_11_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_copy1184_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1185_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1185_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w116_12_c12 :  std_logic;
signal bh86_w117_6_c12 :  std_logic;
signal bh86_w118_8_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_copy1186_c12 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1187_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1187_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w118_9_c12 :  std_logic;
signal bh86_w119_4_c12 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_copy1188_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1189_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1189_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w40_2_c12, bh86_w40_2_c13 :  std_logic;
signal bh86_w41_2_c12, bh86_w41_2_c13 :  std_logic;
signal bh86_w42_2_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_copy1190_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1191_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1191_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w42_3_c12 :  std_logic;
signal bh86_w43_2_c12 :  std_logic;
signal bh86_w44_37_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_copy1192_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1193_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1193_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w44_38_c12 :  std_logic;
signal bh86_w45_33_c12 :  std_logic;
signal bh86_w46_40_c12 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_copy1194_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1195_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1195_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_c12 :  std_logic_vector(2 downto 0);
signal bh86_w46_41_c12 :  std_logic;
signal bh86_w47_44_c12 :  std_logic;
signal bh86_w48_46_c12, bh86_w48_46_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_copy1196_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1197_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1197_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w48_47_c13 :  std_logic;
signal bh86_w49_47_c13 :  std_logic;
signal bh86_w50_46_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_copy1198_c12, Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_copy1198_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1199_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1199_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w50_47_c13 :  std_logic;
signal bh86_w51_42_c13 :  std_logic;
signal bh86_w52_42_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_copy1200_c12, Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_copy1200_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1201_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w51_43_c12, bh86_w51_43_c13 :  std_logic;
signal bh86_w52_43_c12, bh86_w52_43_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_copy1202_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1203_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1203_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w52_44_c13 :  std_logic;
signal bh86_w53_39_c13 :  std_logic;
signal bh86_w54_37_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_copy1204_c12, Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_copy1204_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1205_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w53_40_c12, bh86_w53_40_c13 :  std_logic;
signal bh86_w54_38_c12, bh86_w54_38_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_copy1206_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1207_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1207_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w54_39_c13 :  std_logic;
signal bh86_w55_34_c13 :  std_logic;
signal bh86_w56_29_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_copy1208_c12, Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_copy1208_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1209_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1209_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w55_35_c13 :  std_logic;
signal bh86_w56_30_c13 :  std_logic;
signal bh86_w57_30_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_copy1210_c12, Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_copy1210_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1211_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w56_31_c12, bh86_w56_31_c13 :  std_logic;
signal bh86_w57_31_c12, bh86_w57_31_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_copy1212_c12 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1213_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w57_32_c13 :  std_logic;
signal bh86_w58_23_c13 :  std_logic;
signal bh86_w59_27_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_copy1214_c12, Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_copy1214_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1215_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w58_24_c13 :  std_logic;
signal bh86_w59_28_c13 :  std_logic;
signal bh86_w60_22_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_copy1216_c12, Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_copy1216_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1217_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w59_29_c13 :  std_logic;
signal bh86_w60_23_c13 :  std_logic;
signal bh86_w61_23_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_copy1218_c12, Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_copy1218_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1219_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w60_24_c13 :  std_logic;
signal bh86_w61_24_c13 :  std_logic;
signal bh86_w62_19_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_copy1220_c12, Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_copy1220_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1221_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w61_25_c13 :  std_logic;
signal bh86_w62_20_c13 :  std_logic;
signal bh86_w63_20_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_copy1222_c12, Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_copy1222_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1223_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w62_21_c13 :  std_logic;
signal bh86_w63_21_c13 :  std_logic;
signal bh86_w64_16_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_copy1224_c12, Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_copy1224_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1225_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w63_22_c13 :  std_logic;
signal bh86_w64_17_c13 :  std_logic;
signal bh86_w65_21_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_copy1226_c12, Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_copy1226_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1227_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w64_18_c13 :  std_logic;
signal bh86_w65_22_c13 :  std_logic;
signal bh86_w66_14_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_copy1228_c12, Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_copy1228_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1229_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w65_23_c13 :  std_logic;
signal bh86_w66_15_c13 :  std_logic;
signal bh86_w67_20_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_copy1230_c12, Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_copy1230_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1231_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w66_16_c13 :  std_logic;
signal bh86_w67_21_c13 :  std_logic;
signal bh86_w68_15_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_copy1232_c12, Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_copy1232_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1233_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w67_22_c13 :  std_logic;
signal bh86_w68_16_c13 :  std_logic;
signal bh86_w69_19_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_copy1234_c12, Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_copy1234_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1235_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w68_17_c13 :  std_logic;
signal bh86_w69_20_c13 :  std_logic;
signal bh86_w70_17_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_copy1236_c12, Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_copy1236_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1237_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w69_21_c13 :  std_logic;
signal bh86_w70_18_c13 :  std_logic;
signal bh86_w71_17_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_copy1238_c12, Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_copy1238_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1239_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w70_19_c13 :  std_logic;
signal bh86_w71_18_c13 :  std_logic;
signal bh86_w72_16_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_copy1240_c12, Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_copy1240_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1241_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w71_19_c13 :  std_logic;
signal bh86_w72_17_c13 :  std_logic;
signal bh86_w73_17_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_copy1242_c12, Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_copy1242_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1243_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w72_18_c13 :  std_logic;
signal bh86_w73_18_c13 :  std_logic;
signal bh86_w74_16_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_copy1244_c12, Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_copy1244_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1245_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w73_19_c13 :  std_logic;
signal bh86_w74_17_c13 :  std_logic;
signal bh86_w75_17_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_copy1246_c12, Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_copy1246_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1247_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w74_18_c13 :  std_logic;
signal bh86_w75_18_c13 :  std_logic;
signal bh86_w76_17_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_copy1248_c12, Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_copy1248_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1249_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w75_19_c13 :  std_logic;
signal bh86_w76_18_c13 :  std_logic;
signal bh86_w77_16_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_copy1250_c12, Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_copy1250_c13 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1251_In0_c12 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w76_19_c13 :  std_logic;
signal bh86_w77_17_c13 :  std_logic;
signal bh86_w78_18_c13 :  std_logic;
signal Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_copy1252_c12, Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_copy1252_c13 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1253_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w77_18_c13 :  std_logic;
signal bh86_w78_19_c13 :  std_logic;
signal bh86_w79_16_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_copy1254_c12, Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_copy1254_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1255_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1255_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w78_20_c13 :  std_logic;
signal bh86_w79_17_c13 :  std_logic;
signal bh86_w80_19_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_copy1256_c12, Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_copy1256_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1257_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w79_18_c12, bh86_w79_18_c13 :  std_logic;
signal bh86_w80_20_c12, bh86_w80_20_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_copy1258_c12 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1259_In0_c12 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w80_21_c13 :  std_logic;
signal bh86_w81_15_c13 :  std_logic;
signal bh86_w82_18_c13 :  std_logic;
signal Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_copy1260_c12, Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_copy1260_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1261_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1261_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w81_16_c13 :  std_logic;
signal bh86_w82_19_c13 :  std_logic;
signal bh86_w83_15_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_copy1262_c12, Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_copy1262_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1263_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1263_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w82_20_c13 :  std_logic;
signal bh86_w83_16_c13 :  std_logic;
signal bh86_w84_19_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_copy1264_c12, Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_copy1264_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1265_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w83_17_c12, bh86_w83_17_c13 :  std_logic;
signal bh86_w84_20_c12, bh86_w84_20_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_copy1266_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1267_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1267_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w84_21_c13 :  std_logic;
signal bh86_w85_14_c13 :  std_logic;
signal bh86_w86_18_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_copy1268_c12, Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_copy1268_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1269_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w85_15_c12, bh86_w85_15_c13 :  std_logic;
signal bh86_w86_19_c12, bh86_w86_19_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_copy1270_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1271_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1271_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w86_20_c13 :  std_logic;
signal bh86_w87_16_c13 :  std_logic;
signal bh86_w88_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_copy1272_c12, Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_copy1272_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1273_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_c12 :  std_logic_vector(1 downto 0);
signal bh86_w87_17_c12, bh86_w87_17_c13 :  std_logic;
signal bh86_w88_17_c12, bh86_w88_17_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_copy1274_c12 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1275_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1275_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w88_18_c13 :  std_logic;
signal bh86_w89_15_c13 :  std_logic;
signal bh86_w90_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_copy1276_c12, Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_copy1276_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1277_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w89_16_c13 :  std_logic;
signal bh86_w90_17_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_copy1278_c12, Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_copy1278_c13 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1279_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1279_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w90_18_c13 :  std_logic;
signal bh86_w91_14_c13 :  std_logic;
signal bh86_w92_15_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_copy1280_c12, Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_copy1280_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1281_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1281_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w90_19_c13 :  std_logic;
signal bh86_w91_15_c13 :  std_logic;
signal bh86_w92_16_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_copy1282_c12, Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_copy1282_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1283_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w92_17_c13 :  std_logic;
signal bh86_w93_15_c13 :  std_logic;
signal bh86_w94_14_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_copy1284_c12, Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_copy1284_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1285_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w93_16_c13 :  std_logic;
signal bh86_w94_15_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_copy1286_c12, Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_copy1286_c13 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1287_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c0, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c1, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c2, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c3, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c4, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c5, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c6, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c7, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c8, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c9, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c10, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c11, Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w94_16_c13 :  std_logic;
signal bh86_w95_16_c13 :  std_logic;
signal bh86_w96_14_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_copy1288_c12, Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_copy1288_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1289_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w95_17_c13 :  std_logic;
signal bh86_w96_15_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_copy1290_c12, Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_copy1290_c13 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1291_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w96_16_c13 :  std_logic;
signal bh86_w97_17_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_copy1292_c12, Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_copy1292_c13 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1293_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1293_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w97_18_c13 :  std_logic;
signal bh86_w98_13_c13 :  std_logic;
signal bh86_w99_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_copy1294_c12, Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_copy1294_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1295_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1295_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w99_17_c13 :  std_logic;
signal bh86_w100_13_c13 :  std_logic;
signal bh86_w101_17_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_copy1296_c12, Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_copy1296_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1297_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1297_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w101_18_c13 :  std_logic;
signal bh86_w102_12_c13 :  std_logic;
signal bh86_w103_16_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_copy1298_c12, Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_copy1298_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1299_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1299_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w103_17_c13 :  std_logic;
signal bh86_w104_14_c13 :  std_logic;
signal bh86_w105_14_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_copy1300_c12, Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_copy1300_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1301_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1301_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w105_15_c13 :  std_logic;
signal bh86_w106_13_c13 :  std_logic;
signal bh86_w107_14_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_copy1302_c12, Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_copy1302_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1303_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1303_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w107_15_c13 :  std_logic;
signal bh86_w108_13_c13 :  std_logic;
signal bh86_w109_14_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_copy1304_c12, Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_copy1304_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1305_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1305_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w109_15_c13 :  std_logic;
signal bh86_w110_14_c13 :  std_logic;
signal bh86_w111_13_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_copy1306_c12, Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_copy1306_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1307_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1307_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w111_14_c13 :  std_logic;
signal bh86_w112_15_c13 :  std_logic;
signal bh86_w113_13_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_copy1308_c12, Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_copy1308_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1309_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w113_14_c13 :  std_logic;
signal bh86_w114_16_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_copy1310_c12, Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_copy1310_c13 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1311_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w114_17_c13 :  std_logic;
signal bh86_w115_9_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_copy1312_c12, Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_copy1312_c13 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1313_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1313_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w116_13_c13 :  std_logic;
signal bh86_w117_7_c13 :  std_logic;
signal bh86_w118_10_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_copy1314_c12, Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_copy1314_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1315_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1315_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w118_11_c13 :  std_logic;
signal bh86_w119_5_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_copy1316_c12, Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_copy1316_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1317_In0_c12 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1317_In1_c12 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w42_4_c13 :  std_logic;
signal bh86_w43_3_c13 :  std_logic;
signal bh86_w44_39_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_copy1318_c12, Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_copy1318_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1319_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1319_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w44_40_c13 :  std_logic;
signal bh86_w45_34_c13 :  std_logic;
signal bh86_w46_42_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_copy1320_c12, Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_copy1320_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1321_In0_c12 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1321_In1_c12 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w46_43_c13 :  std_logic;
signal bh86_w47_45_c13 :  std_logic;
signal bh86_w48_48_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_copy1322_c12, Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_copy1322_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1323_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1323_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w48_49_c13 :  std_logic;
signal bh86_w49_48_c13 :  std_logic;
signal bh86_w50_48_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_copy1324_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1325_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1325_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w50_49_c13 :  std_logic;
signal bh86_w51_44_c13 :  std_logic;
signal bh86_w52_45_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_copy1326_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1327_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1327_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w52_46_c13 :  std_logic;
signal bh86_w53_41_c13 :  std_logic;
signal bh86_w54_40_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_copy1328_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1329_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1329_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w54_41_c13 :  std_logic;
signal bh86_w55_36_c13 :  std_logic;
signal bh86_w56_32_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_copy1330_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1331_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c12, Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w56_33_c13 :  std_logic;
signal bh86_w57_33_c13 :  std_logic;
signal bh86_w58_25_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_copy1332_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1333_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1333_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w57_34_c13 :  std_logic;
signal bh86_w58_26_c13 :  std_logic;
signal bh86_w59_30_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_copy1334_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1335_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1335_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w59_31_c13 :  std_logic;
signal bh86_w60_25_c13 :  std_logic;
signal bh86_w61_26_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_copy1336_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1337_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1337_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w61_27_c13 :  std_logic;
signal bh86_w62_22_c13 :  std_logic;
signal bh86_w63_23_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_copy1338_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1339_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1339_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w63_24_c13 :  std_logic;
signal bh86_w64_19_c13 :  std_logic;
signal bh86_w65_24_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_copy1340_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1341_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1341_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w65_25_c13 :  std_logic;
signal bh86_w66_17_c13 :  std_logic;
signal bh86_w67_23_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_copy1342_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1343_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1343_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w67_24_c13 :  std_logic;
signal bh86_w68_18_c13 :  std_logic;
signal bh86_w69_22_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_copy1344_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1345_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1345_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w69_23_c13 :  std_logic;
signal bh86_w70_20_c13 :  std_logic;
signal bh86_w71_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_copy1346_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1347_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1347_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w71_21_c13 :  std_logic;
signal bh86_w72_19_c13 :  std_logic;
signal bh86_w73_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_copy1348_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1349_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1349_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w73_21_c13 :  std_logic;
signal bh86_w74_19_c13 :  std_logic;
signal bh86_w75_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_copy1350_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1351_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1351_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w75_21_c13 :  std_logic;
signal bh86_w76_20_c13 :  std_logic;
signal bh86_w77_19_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_copy1352_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1353_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_c13 :  std_logic_vector(1 downto 0);
signal bh86_w77_20_c13 :  std_logic;
signal bh86_w78_21_c13 :  std_logic;
signal Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_copy1354_c13 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1355_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1355_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w78_22_c13 :  std_logic;
signal bh86_w79_19_c13 :  std_logic;
signal bh86_w80_22_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_copy1356_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1357_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c0, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c1, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c2, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c3, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c4, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c5, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c6, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c7, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c8, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c9, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c10, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c11, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c12, Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w79_20_c13 :  std_logic;
signal bh86_w80_23_c13 :  std_logic;
signal bh86_w81_17_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_copy1358_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1359_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1359_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w80_24_c13 :  std_logic;
signal bh86_w81_18_c13 :  std_logic;
signal bh86_w82_21_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_copy1360_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1361_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1361_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w82_22_c13 :  std_logic;
signal bh86_w83_18_c13 :  std_logic;
signal bh86_w84_22_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_copy1362_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1363_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1363_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w84_23_c13 :  std_logic;
signal bh86_w85_16_c13 :  std_logic;
signal bh86_w86_21_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_copy1364_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1365_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1365_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w86_22_c13 :  std_logic;
signal bh86_w87_18_c13 :  std_logic;
signal bh86_w88_19_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_copy1366_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1367_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1367_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w88_20_c13 :  std_logic;
signal bh86_w89_17_c13 :  std_logic;
signal bh86_w90_20_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_copy1368_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1369_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1369_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w90_21_c13 :  std_logic;
signal bh86_w91_16_c13 :  std_logic;
signal bh86_w92_18_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_copy1370_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1371_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1371_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w92_19_c13 :  std_logic;
signal bh86_w93_17_c13 :  std_logic;
signal bh86_w94_17_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_copy1372_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1373_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1373_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w94_18_c13 :  std_logic;
signal bh86_w95_18_c13 :  std_logic;
signal bh86_w96_17_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_copy1374_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1375_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1375_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w96_18_c13 :  std_logic;
signal bh86_w97_19_c13 :  std_logic;
signal bh86_w98_14_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_copy1376_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1377_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1377_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w98_15_c13 :  std_logic;
signal bh86_w99_18_c13 :  std_logic;
signal bh86_w100_14_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_copy1378_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1379_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1379_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w101_19_c13 :  std_logic;
signal bh86_w102_13_c13 :  std_logic;
signal bh86_w103_18_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_copy1380_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1381_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1381_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w103_19_c13 :  std_logic;
signal bh86_w104_15_c13 :  std_logic;
signal bh86_w105_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_copy1382_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1383_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1383_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w105_17_c13 :  std_logic;
signal bh86_w106_14_c13 :  std_logic;
signal bh86_w107_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_copy1384_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1385_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1385_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w107_17_c13 :  std_logic;
signal bh86_w108_14_c13 :  std_logic;
signal bh86_w109_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_copy1386_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1387_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1387_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w109_17_c13 :  std_logic;
signal bh86_w110_15_c13 :  std_logic;
signal bh86_w111_15_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_copy1388_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1389_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1389_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w111_16_c13 :  std_logic;
signal bh86_w112_16_c13 :  std_logic;
signal bh86_w113_15_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_copy1390_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1391_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1391_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w113_16_c13 :  std_logic;
signal bh86_w114_18_c13 :  std_logic;
signal bh86_w115_10_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_copy1392_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1393_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1393_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w115_11_c13 :  std_logic;
signal bh86_w116_14_c13 :  std_logic;
signal bh86_w117_8_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_copy1394_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1395_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1395_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w118_12_c13 :  std_logic;
signal bh86_w119_6_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_copy1396_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1397_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1397_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w44_41_c13 :  std_logic;
signal bh86_w45_35_c13 :  std_logic;
signal bh86_w46_44_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_copy1398_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1399_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1399_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w46_45_c13 :  std_logic;
signal bh86_w47_46_c13 :  std_logic;
signal bh86_w48_50_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_copy1400_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1401_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1401_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w48_51_c13 :  std_logic;
signal bh86_w49_49_c13 :  std_logic;
signal bh86_w50_50_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_copy1402_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1403_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1403_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w50_51_c13 :  std_logic;
signal bh86_w51_45_c13 :  std_logic;
signal bh86_w52_47_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_copy1404_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1405_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1405_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w52_48_c13 :  std_logic;
signal bh86_w53_42_c13 :  std_logic;
signal bh86_w54_42_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_copy1406_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1407_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1407_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w54_43_c13 :  std_logic;
signal bh86_w55_37_c13 :  std_logic;
signal bh86_w56_34_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_copy1408_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1409_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1409_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w56_35_c13 :  std_logic;
signal bh86_w57_35_c13 :  std_logic;
signal bh86_w58_27_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_copy1410_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1411_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1411_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w58_28_c13 :  std_logic;
signal bh86_w59_32_c13 :  std_logic;
signal bh86_w60_26_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_copy1412_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1413_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1413_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w60_27_c13 :  std_logic;
signal bh86_w61_28_c13 :  std_logic;
signal bh86_w62_23_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_copy1414_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1415_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1415_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w62_24_c13 :  std_logic;
signal bh86_w63_25_c13 :  std_logic;
signal bh86_w64_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_copy1416_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1417_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1417_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w64_21_c13 :  std_logic;
signal bh86_w65_26_c13 :  std_logic;
signal bh86_w66_18_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_copy1418_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1419_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1419_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w66_19_c13 :  std_logic;
signal bh86_w67_25_c13 :  std_logic;
signal bh86_w68_19_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_copy1420_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1421_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1421_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w68_20_c13 :  std_logic;
signal bh86_w69_24_c13 :  std_logic;
signal bh86_w70_21_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_copy1422_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1423_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1423_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w70_22_c13 :  std_logic;
signal bh86_w71_22_c13 :  std_logic;
signal bh86_w72_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_copy1424_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1425_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1425_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w72_21_c13 :  std_logic;
signal bh86_w73_22_c13 :  std_logic;
signal bh86_w74_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_copy1426_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1427_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1427_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w74_21_c13 :  std_logic;
signal bh86_w75_22_c13 :  std_logic;
signal bh86_w76_21_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_copy1428_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1429_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1429_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w76_22_c13 :  std_logic;
signal bh86_w77_21_c13 :  std_logic;
signal bh86_w78_23_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_copy1430_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1431_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1431_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w78_24_c13 :  std_logic;
signal bh86_w79_21_c13 :  std_logic;
signal bh86_w80_25_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_copy1432_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1433_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1433_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w80_26_c13 :  std_logic;
signal bh86_w81_19_c13 :  std_logic;
signal bh86_w82_23_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_copy1434_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1435_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1435_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w82_24_c13 :  std_logic;
signal bh86_w83_19_c13 :  std_logic;
signal bh86_w84_24_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_copy1436_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1437_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1437_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w84_25_c13 :  std_logic;
signal bh86_w85_17_c13 :  std_logic;
signal bh86_w86_23_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_copy1438_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1439_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1439_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w86_24_c13 :  std_logic;
signal bh86_w87_19_c13 :  std_logic;
signal bh86_w88_21_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_copy1440_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1441_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1441_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w88_22_c13 :  std_logic;
signal bh86_w89_18_c13 :  std_logic;
signal bh86_w90_22_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_copy1442_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1443_In0_c13 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1443_In1_c13 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w90_23_c13 :  std_logic;
signal bh86_w91_17_c13 :  std_logic;
signal bh86_w92_20_c13 :  std_logic;
signal Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_copy1444_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1445_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1445_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w92_21_c13 :  std_logic;
signal bh86_w93_18_c13 :  std_logic;
signal bh86_w94_19_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_copy1446_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1447_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1447_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w94_20_c13 :  std_logic;
signal bh86_w95_19_c13 :  std_logic;
signal bh86_w96_19_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_copy1448_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1449_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1449_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w96_20_c13 :  std_logic;
signal bh86_w97_20_c13 :  std_logic;
signal bh86_w98_16_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_copy1450_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1451_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1451_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w98_17_c13 :  std_logic;
signal bh86_w99_19_c13 :  std_logic;
signal bh86_w100_15_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_copy1452_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1453_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1453_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w100_16_c13 :  std_logic;
signal bh86_w101_20_c13 :  std_logic;
signal bh86_w102_14_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_copy1454_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1455_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1455_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w103_20_c13 :  std_logic;
signal bh86_w104_16_c13 :  std_logic;
signal bh86_w105_18_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_copy1456_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1457_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1457_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w105_19_c13 :  std_logic;
signal bh86_w106_15_c13 :  std_logic;
signal bh86_w107_18_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_copy1458_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1459_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1459_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w107_19_c13 :  std_logic;
signal bh86_w108_15_c13 :  std_logic;
signal bh86_w109_18_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_copy1460_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1461_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1461_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w109_19_c13 :  std_logic;
signal bh86_w110_16_c13 :  std_logic;
signal bh86_w111_17_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_copy1462_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1463_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1463_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w111_18_c13 :  std_logic;
signal bh86_w112_17_c13 :  std_logic;
signal bh86_w113_17_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_copy1464_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1465_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1465_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w113_18_c13 :  std_logic;
signal bh86_w114_19_c13 :  std_logic;
signal bh86_w115_12_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_copy1466_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1467_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1467_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w115_13_c13 :  std_logic;
signal bh86_w116_15_c13 :  std_logic;
signal bh86_w117_9_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_copy1468_c13 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1469_In0_c13 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1469_In1_c13 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_c13 :  std_logic_vector(2 downto 0);
signal bh86_w117_10_c13 :  std_logic;
signal bh86_w118_13_c13 :  std_logic;
signal bh86_w119_7_c13 :  std_logic;
signal Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_copy1470_c13 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh86_45_c13, tmp_bitheapResult_bh86_45_c14 :  std_logic_vector(45 downto 0);
signal bitheapFinalAdd_bh86_In0_c13 :  std_logic_vector(74 downto 0);
signal bitheapFinalAdd_bh86_In1_c13 :  std_logic_vector(74 downto 0);
signal bitheapFinalAdd_bh86_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh86_Out_c14 :  std_logic_vector(74 downto 0);
signal bitheapResult_bh86_c14 :  std_logic_vector(119 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh86_w44_30_c1 <= bh86_w44_30_c0;
               bh86_w46_20_c1 <= bh86_w46_20_c0;
               bh86_w47_24_c1 <= bh86_w47_24_c0;
               bh86_w49_22_c1 <= bh86_w49_22_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c0;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c1 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c0;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c1 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c0;
            end if;
            if ce_2 = '1' then
               bh86_w44_30_c2 <= bh86_w44_30_c1;
               bh86_w46_20_c2 <= bh86_w46_20_c1;
               bh86_w47_24_c2 <= bh86_w47_24_c1;
               bh86_w49_22_c2 <= bh86_w49_22_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c1;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c2 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c1;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c2 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c1;
            end if;
            if ce_3 = '1' then
               bh86_w44_30_c3 <= bh86_w44_30_c2;
               bh86_w46_20_c3 <= bh86_w46_20_c2;
               bh86_w47_24_c3 <= bh86_w47_24_c2;
               bh86_w49_22_c3 <= bh86_w49_22_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c2;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c3 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c2;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c3 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c2;
            end if;
            if ce_4 = '1' then
               bh86_w44_30_c4 <= bh86_w44_30_c3;
               bh86_w46_20_c4 <= bh86_w46_20_c3;
               bh86_w47_24_c4 <= bh86_w47_24_c3;
               bh86_w49_22_c4 <= bh86_w49_22_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c3;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c4 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c3;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c4 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c3;
            end if;
            if ce_5 = '1' then
               bh86_w44_30_c5 <= bh86_w44_30_c4;
               bh86_w46_20_c5 <= bh86_w46_20_c4;
               bh86_w47_24_c5 <= bh86_w47_24_c4;
               bh86_w49_22_c5 <= bh86_w49_22_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c4;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c5 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c4;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c5 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c4;
            end if;
            if ce_6 = '1' then
               bh86_w44_30_c6 <= bh86_w44_30_c5;
               bh86_w46_20_c6 <= bh86_w46_20_c5;
               bh86_w47_24_c6 <= bh86_w47_24_c5;
               bh86_w49_22_c6 <= bh86_w49_22_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c5;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c6 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c5;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c6 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c5;
            end if;
            if ce_7 = '1' then
               bh86_w44_30_c7 <= bh86_w44_30_c6;
               bh86_w46_20_c7 <= bh86_w46_20_c6;
               bh86_w47_24_c7 <= bh86_w47_24_c6;
               bh86_w49_22_c7 <= bh86_w49_22_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c6;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c7 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c6;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c7 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c6;
            end if;
            if ce_8 = '1' then
               bh86_w44_30_c8 <= bh86_w44_30_c7;
               bh86_w46_20_c8 <= bh86_w46_20_c7;
               bh86_w47_24_c8 <= bh86_w47_24_c7;
               bh86_w49_22_c8 <= bh86_w49_22_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c7;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c8 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c7;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c8 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c7;
            end if;
            if ce_9 = '1' then
               bh86_w44_30_c9 <= bh86_w44_30_c8;
               bh86_w46_20_c9 <= bh86_w46_20_c8;
               bh86_w47_24_c9 <= bh86_w47_24_c8;
               bh86_w49_22_c9 <= bh86_w49_22_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c8;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c9 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c8;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c9 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c8;
            end if;
            if ce_10 = '1' then
               bh86_w44_30_c10 <= bh86_w44_30_c9;
               bh86_w46_20_c10 <= bh86_w46_20_c9;
               bh86_w47_24_c10 <= bh86_w47_24_c9;
               bh86_w49_22_c10 <= bh86_w49_22_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c9;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c10 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c9;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c10 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c9;
            end if;
            if ce_11 = '1' then
               bh86_w44_30_c11 <= bh86_w44_30_c10;
               bh86_w46_20_c11 <= bh86_w46_20_c10;
               bh86_w47_24_c11 <= bh86_w47_24_c10;
               bh86_w49_22_c11 <= bh86_w49_22_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c10;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c11 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c10;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c11 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c10;
            end if;
            if ce_12 = '1' then
               bh86_w44_12_c12 <= bh86_w44_12_c11;
               bh86_w46_7_c12 <= bh86_w46_7_c11;
               bh86_w52_13_c12 <= bh86_w52_13_c11;
               bh86_w104_5_c12 <= bh86_w104_5_c11;
               bh86_w115_2_c12 <= bh86_w115_2_c11;
               bh86_w118_0_c12 <= bh86_w118_0_c11;
               bh86_w87_7_c12 <= bh86_w87_7_c11;
               bh86_w101_5_c12 <= bh86_w101_5_c11;
               bh86_w70_8_c12 <= bh86_w70_8_c11;
               bh86_w84_7_c12 <= bh86_w84_7_c11;
               bh86_w58_11_c12 <= bh86_w58_11_c11;
               bh86_w63_8_c12 <= bh86_w63_8_c11;
               bh86_w65_8_c12 <= bh86_w65_8_c11;
               bh86_w67_8_c12 <= bh86_w67_8_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_copy618_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_copy618_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_copy620_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_copy620_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_copy622_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_copy622_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_copy624_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_copy624_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_copy628_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_copy628_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_copy630_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_copy630_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_copy632_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_copy632_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_copy634_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_copy634_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_copy636_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_copy636_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_copy638_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_copy638_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_copy640_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_copy640_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_copy642_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_copy642_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_copy644_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_copy644_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_copy646_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_copy646_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_copy648_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_copy648_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_copy652_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_copy652_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_copy654_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_copy654_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_copy656_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_copy656_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_copy658_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_copy658_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_copy660_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_copy660_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_copy662_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_copy662_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_copy664_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_copy664_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_copy666_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_copy666_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_copy668_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_copy668_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_copy670_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_copy670_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_copy672_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_copy672_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_copy674_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_copy674_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_copy676_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_copy676_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_copy678_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_copy678_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_copy680_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_copy680_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_copy682_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_copy682_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_copy684_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_copy684_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_copy686_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_copy686_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_copy688_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_copy688_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_copy690_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_copy690_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_copy692_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_copy692_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_copy694_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_copy694_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_copy696_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_copy696_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_copy698_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_copy698_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_copy700_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_copy700_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_copy702_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_copy702_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_copy704_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_copy704_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_copy706_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_copy706_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_copy708_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_copy708_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_copy710_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_copy710_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_copy714_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_copy714_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_copy716_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_copy716_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_copy718_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_copy718_c11;
               Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_copy720_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_copy720_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_copy722_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_copy722_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_copy724_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_copy724_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_copy726_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_copy726_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_copy728_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_copy728_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_copy730_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_copy730_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_copy732_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_copy732_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_copy734_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_copy734_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_copy736_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_copy736_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_copy738_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_copy738_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_copy740_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_copy740_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_copy742_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_copy742_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_copy744_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_copy744_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_copy746_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_copy746_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_copy748_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_copy748_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_copy750_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_copy750_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_copy752_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_copy752_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_copy754_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_copy754_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_copy756_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_copy756_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_copy758_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_copy758_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_copy760_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_copy760_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_copy762_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_copy762_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_copy764_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_copy764_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_copy766_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_copy766_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_copy768_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_copy768_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_copy770_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_copy770_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_copy772_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_copy772_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_copy774_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_copy774_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_copy776_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_copy776_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_copy778_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_copy778_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_copy780_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_copy780_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_copy782_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_copy782_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_copy784_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_copy784_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_copy786_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_copy786_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_copy788_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_copy788_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_copy790_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_copy790_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_copy792_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_copy792_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_copy794_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_copy794_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_copy796_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_copy796_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_copy798_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_copy798_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_copy800_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_copy800_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_copy802_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_copy802_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_copy804_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_copy804_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_copy806_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_copy806_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_copy808_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_copy808_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_copy810_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_copy810_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_copy812_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_copy812_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_copy814_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_copy814_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_copy816_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_copy816_c11;
               Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_copy818_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_copy818_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_copy820_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_copy820_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_copy822_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_copy822_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_copy824_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_copy824_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_copy826_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_copy826_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid875_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid875_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid953_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid953_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c11;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c11;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c11;
            end if;
            if ce_13 = '1' then
               bh86_w33_0_c13 <= bh86_w33_0_c12;
               bh86_w34_0_c13 <= bh86_w34_0_c12;
               bh86_w35_0_c13 <= bh86_w35_0_c12;
               bh86_w36_0_c13 <= bh86_w36_0_c12;
               bh86_w37_0_c13 <= bh86_w37_0_c12;
               bh86_w38_0_c13 <= bh86_w38_0_c12;
               bh86_w39_0_c13 <= bh86_w39_0_c12;
               bh86_w49_0_c13 <= bh86_w49_0_c12;
               bh86_w50_1_c13 <= bh86_w50_1_c12;
               bh86_w52_1_c13 <= bh86_w52_1_c12;
               bh86_w54_1_c13 <= bh86_w54_1_c12;
               bh86_w98_0_c13 <= bh86_w98_0_c12;
               bh86_w84_2_c13 <= bh86_w84_2_c12;
               bh86_w86_2_c13 <= bh86_w86_2_c12;
               bh86_w78_3_c13 <= bh86_w78_3_c12;
               bh86_w79_3_c13 <= bh86_w79_3_c12;
               bh86_w88_15_c13 <= bh86_w88_15_c12;
               bh86_w115_8_c13 <= bh86_w115_8_c12;
               bh86_w40_2_c13 <= bh86_w40_2_c12;
               bh86_w41_2_c13 <= bh86_w41_2_c12;
               bh86_w48_46_c13 <= bh86_w48_46_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_copy1198_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_copy1198_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_copy1200_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_copy1200_c12;
               bh86_w51_43_c13 <= bh86_w51_43_c12;
               bh86_w52_43_c13 <= bh86_w52_43_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_copy1204_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_copy1204_c12;
               bh86_w53_40_c13 <= bh86_w53_40_c12;
               bh86_w54_38_c13 <= bh86_w54_38_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_copy1208_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_copy1208_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_copy1210_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_copy1210_c12;
               bh86_w56_31_c13 <= bh86_w56_31_c12;
               bh86_w57_31_c13 <= bh86_w57_31_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_copy1214_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_copy1214_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_copy1216_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_copy1216_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_copy1218_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_copy1218_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_copy1220_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_copy1220_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_copy1222_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_copy1222_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_copy1224_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_copy1224_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_copy1226_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_copy1226_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_copy1228_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_copy1228_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_copy1230_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_copy1230_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_copy1232_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_copy1232_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_copy1234_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_copy1234_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_copy1236_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_copy1236_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_copy1238_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_copy1238_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_copy1240_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_copy1240_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_copy1242_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_copy1242_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_copy1244_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_copy1244_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_copy1246_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_copy1246_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_copy1248_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_copy1248_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_copy1250_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_copy1250_c12;
               Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_copy1252_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_copy1252_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_copy1254_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_copy1254_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_copy1256_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_copy1256_c12;
               bh86_w79_18_c13 <= bh86_w79_18_c12;
               bh86_w80_20_c13 <= bh86_w80_20_c12;
               Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_copy1260_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_copy1260_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_copy1262_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_copy1262_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_copy1264_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_copy1264_c12;
               bh86_w83_17_c13 <= bh86_w83_17_c12;
               bh86_w84_20_c13 <= bh86_w84_20_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_copy1268_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_copy1268_c12;
               bh86_w85_15_c13 <= bh86_w85_15_c12;
               bh86_w86_19_c13 <= bh86_w86_19_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_copy1272_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_copy1272_c12;
               bh86_w87_17_c13 <= bh86_w87_17_c12;
               bh86_w88_17_c13 <= bh86_w88_17_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_copy1276_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_copy1276_c12;
               Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_copy1278_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_copy1278_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_copy1280_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_copy1280_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_copy1282_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_copy1282_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_copy1284_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_copy1284_c12;
               Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_copy1286_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_copy1286_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_copy1288_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_copy1288_c12;
               Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_copy1290_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_copy1290_c12;
               Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_copy1292_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_copy1292_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_copy1294_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_copy1294_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_copy1296_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_copy1296_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_copy1298_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_copy1298_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_copy1300_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_copy1300_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_copy1302_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_copy1302_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_copy1304_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_copy1304_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_copy1306_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_copy1306_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_copy1308_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_copy1308_c12;
               Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_copy1310_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_copy1310_c12;
               Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_copy1312_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_copy1312_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_copy1314_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_copy1314_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_copy1316_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_copy1316_c12;
               Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_copy1318_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_copy1318_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_copy1320_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_copy1320_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_copy1322_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_copy1322_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c12;
               Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c12;
            end if;
            if ce_14 = '1' then
               tmp_bitheapResult_bh86_45_c14 <= tmp_bitheapResult_bh86_45_c13;
            end if;
         end if;
      end process;
   XX_m85_c11 <= X ;
   YY_m85_c0 <= Y ;
   tile_0_X_c11 <= X(66 downto 50);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid88
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 X => tile_0_X_c11,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c12);

   tile_0_filtered_output_c12 <= unsigned(tile_0_output_c12(40 downto 0));
   bh86_w50_0_c12 <= tile_0_filtered_output_c12(0);
   bh86_w51_0_c12 <= tile_0_filtered_output_c12(1);
   bh86_w52_0_c12 <= tile_0_filtered_output_c12(2);
   bh86_w53_0_c12 <= tile_0_filtered_output_c12(3);
   bh86_w54_0_c12 <= tile_0_filtered_output_c12(4);
   bh86_w55_0_c12 <= tile_0_filtered_output_c12(5);
   bh86_w56_0_c12 <= tile_0_filtered_output_c12(6);
   bh86_w57_0_c12 <= tile_0_filtered_output_c12(7);
   bh86_w58_0_c12 <= tile_0_filtered_output_c12(8);
   bh86_w59_0_c12 <= tile_0_filtered_output_c12(9);
   bh86_w60_0_c12 <= tile_0_filtered_output_c12(10);
   bh86_w61_0_c12 <= tile_0_filtered_output_c12(11);
   bh86_w62_0_c12 <= tile_0_filtered_output_c12(12);
   bh86_w63_0_c12 <= tile_0_filtered_output_c12(13);
   bh86_w64_0_c12 <= tile_0_filtered_output_c12(14);
   bh86_w65_0_c12 <= tile_0_filtered_output_c12(15);
   bh86_w66_0_c12 <= tile_0_filtered_output_c12(16);
   bh86_w67_0_c12 <= tile_0_filtered_output_c12(17);
   bh86_w68_0_c12 <= tile_0_filtered_output_c12(18);
   bh86_w69_0_c12 <= tile_0_filtered_output_c12(19);
   bh86_w70_0_c12 <= tile_0_filtered_output_c12(20);
   bh86_w71_0_c12 <= tile_0_filtered_output_c12(21);
   bh86_w72_0_c12 <= tile_0_filtered_output_c12(22);
   bh86_w73_0_c12 <= tile_0_filtered_output_c12(23);
   bh86_w74_0_c12 <= tile_0_filtered_output_c12(24);
   bh86_w75_0_c12 <= tile_0_filtered_output_c12(25);
   bh86_w76_0_c12 <= tile_0_filtered_output_c12(26);
   bh86_w77_0_c12 <= tile_0_filtered_output_c12(27);
   bh86_w78_0_c12 <= tile_0_filtered_output_c12(28);
   bh86_w79_0_c12 <= tile_0_filtered_output_c12(29);
   bh86_w80_0_c12 <= tile_0_filtered_output_c12(30);
   bh86_w81_0_c12 <= tile_0_filtered_output_c12(31);
   bh86_w82_0_c12 <= tile_0_filtered_output_c12(32);
   bh86_w83_0_c12 <= tile_0_filtered_output_c12(33);
   bh86_w84_0_c12 <= tile_0_filtered_output_c12(34);
   bh86_w85_0_c12 <= tile_0_filtered_output_c12(35);
   bh86_w86_0_c12 <= tile_0_filtered_output_c12(36);
   bh86_w87_0_c12 <= tile_0_filtered_output_c12(37);
   bh86_w88_0_c12 <= tile_0_filtered_output_c12(38);
   bh86_w89_0_c12 <= tile_0_filtered_output_c12(39);
   bh86_w90_0_c12 <= tile_0_filtered_output_c12(40);
   tile_1_X_c11 <= X(49 downto 33);
   tile_1_Y_c0 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_Freq300_uid90
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 X => tile_1_X_c11,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c12);

   tile_1_filtered_output_c12 <= unsigned(tile_1_output_c12(40 downto 0));
   bh86_w33_0_c12 <= tile_1_filtered_output_c12(0);
   bh86_w34_0_c12 <= tile_1_filtered_output_c12(1);
   bh86_w35_0_c12 <= tile_1_filtered_output_c12(2);
   bh86_w36_0_c12 <= tile_1_filtered_output_c12(3);
   bh86_w37_0_c12 <= tile_1_filtered_output_c12(4);
   bh86_w38_0_c12 <= tile_1_filtered_output_c12(5);
   bh86_w39_0_c12 <= tile_1_filtered_output_c12(6);
   bh86_w40_0_c12 <= tile_1_filtered_output_c12(7);
   bh86_w41_0_c12 <= tile_1_filtered_output_c12(8);
   bh86_w42_0_c12 <= tile_1_filtered_output_c12(9);
   bh86_w43_0_c12 <= tile_1_filtered_output_c12(10);
   bh86_w44_0_c12 <= tile_1_filtered_output_c12(11);
   bh86_w45_0_c12 <= tile_1_filtered_output_c12(12);
   bh86_w46_0_c12 <= tile_1_filtered_output_c12(13);
   bh86_w47_0_c12 <= tile_1_filtered_output_c12(14);
   bh86_w48_0_c12 <= tile_1_filtered_output_c12(15);
   bh86_w49_0_c12 <= tile_1_filtered_output_c12(16);
   bh86_w50_1_c12 <= tile_1_filtered_output_c12(17);
   bh86_w51_1_c12 <= tile_1_filtered_output_c12(18);
   bh86_w52_1_c12 <= tile_1_filtered_output_c12(19);
   bh86_w53_1_c12 <= tile_1_filtered_output_c12(20);
   bh86_w54_1_c12 <= tile_1_filtered_output_c12(21);
   bh86_w55_1_c12 <= tile_1_filtered_output_c12(22);
   bh86_w56_1_c12 <= tile_1_filtered_output_c12(23);
   bh86_w57_1_c12 <= tile_1_filtered_output_c12(24);
   bh86_w58_1_c12 <= tile_1_filtered_output_c12(25);
   bh86_w59_1_c12 <= tile_1_filtered_output_c12(26);
   bh86_w60_1_c12 <= tile_1_filtered_output_c12(27);
   bh86_w61_1_c12 <= tile_1_filtered_output_c12(28);
   bh86_w62_1_c12 <= tile_1_filtered_output_c12(29);
   bh86_w63_1_c12 <= tile_1_filtered_output_c12(30);
   bh86_w64_1_c12 <= tile_1_filtered_output_c12(31);
   bh86_w65_1_c12 <= tile_1_filtered_output_c12(32);
   bh86_w66_1_c12 <= tile_1_filtered_output_c12(33);
   bh86_w67_1_c12 <= tile_1_filtered_output_c12(34);
   bh86_w68_1_c12 <= tile_1_filtered_output_c12(35);
   bh86_w69_1_c12 <= tile_1_filtered_output_c12(36);
   bh86_w70_1_c12 <= tile_1_filtered_output_c12(37);
   bh86_w71_1_c12 <= tile_1_filtered_output_c12(38);
   bh86_w72_1_c12 <= tile_1_filtered_output_c12(39);
   bh86_w73_1_c12 <= tile_1_filtered_output_c12(40);
   tile_2_X_c11 <= X(32 downto 32);
   tile_2_Y_c0 <= Y(12 downto 12);
   tile_2_mult: IntMultiplierLUT_1x1_Freq300_uid92
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_2_X_c11,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c11);

   tile_2_filtered_output_c11 <= unsigned(tile_2_output_c11(0 downto 0));
   bh86_w44_1_c11 <= tile_2_filtered_output_c11(0);
   tile_3_X_c11 <= X(32 downto 31);
   tile_3_Y_c0 <= Y(13 downto 13);
   tile_3_mult: IntMultiplierLUT_2x1_Freq300_uid94
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_3_X_c11,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c11);

   tile_3_filtered_output_c11 <= unsigned(tile_3_output_c11(1 downto 0));
   bh86_w44_2_c11 <= tile_3_filtered_output_c11(0);
   bh86_w45_1_c11 <= tile_3_filtered_output_c11(1);
   tile_4_X_c11 <= X(29 downto 29);
   tile_4_Y_c0 <= Y(15 downto 15);
   tile_4_mult: IntMultiplierLUT_1x1_Freq300_uid96
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_4_X_c11,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c11);

   tile_4_filtered_output_c11 <= unsigned(tile_4_output_c11(0 downto 0));
   bh86_w44_3_c11 <= tile_4_filtered_output_c11(0);
   tile_5_X_c11 <= X(32 downto 30);
   tile_5_Y_c0 <= Y(15 downto 14);
   tile_5_mult: IntMultiplierLUT_3x2_Freq300_uid98
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_5_X_c11,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c11);

   tile_5_filtered_output_c11 <= unsigned(tile_5_output_c11(4 downto 0));
   bh86_w44_4_c11 <= tile_5_filtered_output_c11(0);
   bh86_w45_2_c11 <= tile_5_filtered_output_c11(1);
   bh86_w46_1_c11 <= tile_5_filtered_output_c11(2);
   bh86_w47_1_c11 <= tile_5_filtered_output_c11(3);
   bh86_w48_1_c11 <= tile_5_filtered_output_c11(4);
   tile_6_X_c11 <= X(27 downto 27);
   tile_6_Y_c0 <= Y(17 downto 17);
   tile_6_mult: IntMultiplierLUT_1x1_Freq300_uid103
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_6_X_c11,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c11);

   tile_6_filtered_output_c11 <= unsigned(tile_6_output_c11(0 downto 0));
   bh86_w44_5_c11 <= tile_6_filtered_output_c11(0);
   tile_7_X_c11 <= X(29 downto 28);
   tile_7_Y_c0 <= Y(17 downto 16);
   tile_7_mult: IntMultiplierLUT_2x2_Freq300_uid105
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_7_X_c11,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c11);

   tile_7_filtered_output_c11 <= unsigned(tile_7_output_c11(3 downto 0));
   bh86_w44_6_c11 <= tile_7_filtered_output_c11(0);
   bh86_w45_3_c11 <= tile_7_filtered_output_c11(1);
   bh86_w46_2_c11 <= tile_7_filtered_output_c11(2);
   bh86_w47_2_c11 <= tile_7_filtered_output_c11(3);
   tile_8_X_c11 <= X(32 downto 30);
   tile_8_Y_c0 <= Y(17 downto 16);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid110
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_8_X_c11,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c11);

   tile_8_filtered_output_c11 <= unsigned(tile_8_output_c11(4 downto 0));
   bh86_w46_3_c11 <= tile_8_filtered_output_c11(0);
   bh86_w47_3_c11 <= tile_8_filtered_output_c11(1);
   bh86_w48_2_c11 <= tile_8_filtered_output_c11(2);
   bh86_w49_1_c11 <= tile_8_filtered_output_c11(3);
   bh86_w50_2_c11 <= tile_8_filtered_output_c11(4);
   tile_9_X_c11 <= X(26 downto 26);
   tile_9_Y_c0 <= Y(18 downto 18);
   tile_9_mult: IntMultiplierLUT_1x1_Freq300_uid115
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_9_X_c11,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c11);

   tile_9_filtered_output_c11 <= unsigned(tile_9_output_c11(0 downto 0));
   bh86_w44_7_c11 <= tile_9_filtered_output_c11(0);
   tile_10_X_c11 <= X(26 downto 25);
   tile_10_Y_c0 <= Y(19 downto 19);
   tile_10_mult: IntMultiplierLUT_2x1_Freq300_uid117
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_10_X_c11,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c11);

   tile_10_filtered_output_c11 <= unsigned(tile_10_output_c11(1 downto 0));
   bh86_w44_8_c11 <= tile_10_filtered_output_c11(0);
   bh86_w45_4_c11 <= tile_10_filtered_output_c11(1);
   tile_11_X_c11 <= X(29 downto 27);
   tile_11_Y_c0 <= Y(19 downto 18);
   tile_11_mult: IntMultiplierLUT_3x2_Freq300_uid119
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_11_X_c11,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c11);

   tile_11_filtered_output_c11 <= unsigned(tile_11_output_c11(4 downto 0));
   bh86_w45_5_c11 <= tile_11_filtered_output_c11(0);
   bh86_w46_4_c11 <= tile_11_filtered_output_c11(1);
   bh86_w47_4_c11 <= tile_11_filtered_output_c11(2);
   bh86_w48_3_c11 <= tile_11_filtered_output_c11(3);
   bh86_w49_2_c11 <= tile_11_filtered_output_c11(4);
   tile_12_X_c11 <= X(32 downto 30);
   tile_12_Y_c0 <= Y(19 downto 18);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid124
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_12_X_c11,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c11);

   tile_12_filtered_output_c11 <= unsigned(tile_12_output_c11(4 downto 0));
   bh86_w48_4_c11 <= tile_12_filtered_output_c11(0);
   bh86_w49_3_c11 <= tile_12_filtered_output_c11(1);
   bh86_w50_3_c11 <= tile_12_filtered_output_c11(2);
   bh86_w51_2_c11 <= tile_12_filtered_output_c11(3);
   bh86_w52_2_c11 <= tile_12_filtered_output_c11(4);
   tile_13_X_c11 <= X(23 downto 23);
   tile_13_Y_c0 <= Y(21 downto 21);
   tile_13_mult: IntMultiplierLUT_1x1_Freq300_uid129
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_13_X_c11,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c11);

   tile_13_filtered_output_c11 <= unsigned(tile_13_output_c11(0 downto 0));
   bh86_w44_9_c11 <= tile_13_filtered_output_c11(0);
   tile_14_X_c11 <= X(26 downto 24);
   tile_14_Y_c0 <= Y(21 downto 20);
   tile_14_mult: IntMultiplierLUT_3x2_Freq300_uid131
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_14_X_c11,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c11);

   tile_14_filtered_output_c11 <= unsigned(tile_14_output_c11(4 downto 0));
   bh86_w44_10_c11 <= tile_14_filtered_output_c11(0);
   bh86_w45_6_c11 <= tile_14_filtered_output_c11(1);
   bh86_w46_5_c11 <= tile_14_filtered_output_c11(2);
   bh86_w47_5_c11 <= tile_14_filtered_output_c11(3);
   bh86_w48_5_c11 <= tile_14_filtered_output_c11(4);
   tile_15_X_c11 <= X(29 downto 27);
   tile_15_Y_c0 <= Y(21 downto 20);
   tile_15_mult: IntMultiplierLUT_3x2_Freq300_uid136
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_15_X_c11,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c11);

   tile_15_filtered_output_c11 <= unsigned(tile_15_output_c11(4 downto 0));
   bh86_w47_6_c11 <= tile_15_filtered_output_c11(0);
   bh86_w48_6_c11 <= tile_15_filtered_output_c11(1);
   bh86_w49_4_c11 <= tile_15_filtered_output_c11(2);
   bh86_w50_4_c11 <= tile_15_filtered_output_c11(3);
   bh86_w51_3_c11 <= tile_15_filtered_output_c11(4);
   tile_16_X_c11 <= X(32 downto 30);
   tile_16_Y_c0 <= Y(21 downto 20);
   tile_16_mult: IntMultiplierLUT_3x2_Freq300_uid141
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_16_X_c11,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c11);

   tile_16_filtered_output_c11 <= unsigned(tile_16_output_c11(4 downto 0));
   bh86_w50_5_c11 <= tile_16_filtered_output_c11(0);
   bh86_w51_4_c11 <= tile_16_filtered_output_c11(1);
   bh86_w52_3_c11 <= tile_16_filtered_output_c11(2);
   bh86_w53_2_c11 <= tile_16_filtered_output_c11(3);
   bh86_w54_2_c11 <= tile_16_filtered_output_c11(4);
   tile_17_X_c11 <= X(21 downto 21);
   tile_17_Y_c0 <= Y(23 downto 23);
   tile_17_mult: IntMultiplierLUT_1x1_Freq300_uid146
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_17_X_c11,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c11);

   tile_17_filtered_output_c11 <= unsigned(tile_17_output_c11(0 downto 0));
   bh86_w44_11_c11 <= tile_17_filtered_output_c11(0);
   tile_18_X_c11 <= X(23 downto 22);
   tile_18_Y_c0 <= Y(23 downto 22);
   tile_18_mult: IntMultiplierLUT_2x2_Freq300_uid148
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_18_X_c11,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c11);

   tile_18_filtered_output_c11 <= unsigned(tile_18_output_c11(3 downto 0));
   bh86_w44_12_c11 <= tile_18_filtered_output_c11(0);
   bh86_w45_7_c11 <= tile_18_filtered_output_c11(1);
   bh86_w46_6_c11 <= tile_18_filtered_output_c11(2);
   bh86_w47_7_c11 <= tile_18_filtered_output_c11(3);
   tile_19_X_c11 <= X(26 downto 24);
   tile_19_Y_c0 <= Y(23 downto 22);
   tile_19_mult: IntMultiplierLUT_3x2_Freq300_uid153
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_19_X_c11,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c11);

   tile_19_filtered_output_c11 <= unsigned(tile_19_output_c11(4 downto 0));
   bh86_w46_7_c11 <= tile_19_filtered_output_c11(0);
   bh86_w47_8_c11 <= tile_19_filtered_output_c11(1);
   bh86_w48_7_c11 <= tile_19_filtered_output_c11(2);
   bh86_w49_5_c11 <= tile_19_filtered_output_c11(3);
   bh86_w50_6_c11 <= tile_19_filtered_output_c11(4);
   tile_20_X_c11 <= X(29 downto 27);
   tile_20_Y_c0 <= Y(23 downto 22);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid158
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_20_X_c11,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c11);

   tile_20_filtered_output_c11 <= unsigned(tile_20_output_c11(4 downto 0));
   bh86_w49_6_c11 <= tile_20_filtered_output_c11(0);
   bh86_w50_7_c11 <= tile_20_filtered_output_c11(1);
   bh86_w51_5_c11 <= tile_20_filtered_output_c11(2);
   bh86_w52_4_c11 <= tile_20_filtered_output_c11(3);
   bh86_w53_3_c11 <= tile_20_filtered_output_c11(4);
   tile_21_X_c11 <= X(32 downto 30);
   tile_21_Y_c0 <= Y(23 downto 22);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid163
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_21_X_c11,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c11);

   tile_21_filtered_output_c11 <= unsigned(tile_21_output_c11(4 downto 0));
   bh86_w52_5_c11 <= tile_21_filtered_output_c11(0);
   bh86_w53_4_c11 <= tile_21_filtered_output_c11(1);
   bh86_w54_3_c11 <= tile_21_filtered_output_c11(2);
   bh86_w55_2_c11 <= tile_21_filtered_output_c11(3);
   bh86_w56_2_c11 <= tile_21_filtered_output_c11(4);
   tile_22_X_c11 <= X(66 downto 50);
   tile_22_Y_c0 <= Y(47 downto 24);
   tile_22_mult: DSPBlock_17x24_Freq300_uid168
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 X => tile_22_X_c11,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c12);

   tile_22_filtered_output_c12 <= unsigned(tile_22_output_c12(40 downto 0));
   bh86_w74_1_c12 <= tile_22_filtered_output_c12(0);
   bh86_w75_1_c12 <= tile_22_filtered_output_c12(1);
   bh86_w76_1_c12 <= tile_22_filtered_output_c12(2);
   bh86_w77_1_c12 <= tile_22_filtered_output_c12(3);
   bh86_w78_1_c12 <= tile_22_filtered_output_c12(4);
   bh86_w79_1_c12 <= tile_22_filtered_output_c12(5);
   bh86_w80_1_c12 <= tile_22_filtered_output_c12(6);
   bh86_w81_1_c12 <= tile_22_filtered_output_c12(7);
   bh86_w82_1_c12 <= tile_22_filtered_output_c12(8);
   bh86_w83_1_c12 <= tile_22_filtered_output_c12(9);
   bh86_w84_1_c12 <= tile_22_filtered_output_c12(10);
   bh86_w85_1_c12 <= tile_22_filtered_output_c12(11);
   bh86_w86_1_c12 <= tile_22_filtered_output_c12(12);
   bh86_w87_1_c12 <= tile_22_filtered_output_c12(13);
   bh86_w88_1_c12 <= tile_22_filtered_output_c12(14);
   bh86_w89_1_c12 <= tile_22_filtered_output_c12(15);
   bh86_w90_1_c12 <= tile_22_filtered_output_c12(16);
   bh86_w91_0_c12 <= tile_22_filtered_output_c12(17);
   bh86_w92_0_c12 <= tile_22_filtered_output_c12(18);
   bh86_w93_0_c12 <= tile_22_filtered_output_c12(19);
   bh86_w94_0_c12 <= tile_22_filtered_output_c12(20);
   bh86_w95_0_c12 <= tile_22_filtered_output_c12(21);
   bh86_w96_0_c12 <= tile_22_filtered_output_c12(22);
   bh86_w97_0_c12 <= tile_22_filtered_output_c12(23);
   bh86_w98_0_c12 <= tile_22_filtered_output_c12(24);
   bh86_w99_0_c12 <= tile_22_filtered_output_c12(25);
   bh86_w100_0_c12 <= tile_22_filtered_output_c12(26);
   bh86_w101_0_c12 <= tile_22_filtered_output_c12(27);
   bh86_w102_0_c12 <= tile_22_filtered_output_c12(28);
   bh86_w103_0_c12 <= tile_22_filtered_output_c12(29);
   bh86_w104_0_c12 <= tile_22_filtered_output_c12(30);
   bh86_w105_0_c12 <= tile_22_filtered_output_c12(31);
   bh86_w106_0_c12 <= tile_22_filtered_output_c12(32);
   bh86_w107_0_c12 <= tile_22_filtered_output_c12(33);
   bh86_w108_0_c12 <= tile_22_filtered_output_c12(34);
   bh86_w109_0_c12 <= tile_22_filtered_output_c12(35);
   bh86_w110_0_c12 <= tile_22_filtered_output_c12(36);
   bh86_w111_0_c12 <= tile_22_filtered_output_c12(37);
   bh86_w112_0_c12 <= tile_22_filtered_output_c12(38);
   bh86_w113_0_c12 <= tile_22_filtered_output_c12(39);
   bh86_w114_0_c12 <= tile_22_filtered_output_c12(40);
   tile_23_X_c11 <= X(49 downto 33);
   tile_23_Y_c0 <= Y(47 downto 24);
   tile_23_mult: DSPBlock_17x24_Freq300_uid170
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 X => tile_23_X_c11,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c12);

   tile_23_filtered_output_c12 <= unsigned(tile_23_output_c12(40 downto 0));
   bh86_w57_2_c12 <= tile_23_filtered_output_c12(0);
   bh86_w58_2_c12 <= tile_23_filtered_output_c12(1);
   bh86_w59_2_c12 <= tile_23_filtered_output_c12(2);
   bh86_w60_2_c12 <= tile_23_filtered_output_c12(3);
   bh86_w61_2_c12 <= tile_23_filtered_output_c12(4);
   bh86_w62_2_c12 <= tile_23_filtered_output_c12(5);
   bh86_w63_2_c12 <= tile_23_filtered_output_c12(6);
   bh86_w64_2_c12 <= tile_23_filtered_output_c12(7);
   bh86_w65_2_c12 <= tile_23_filtered_output_c12(8);
   bh86_w66_2_c12 <= tile_23_filtered_output_c12(9);
   bh86_w67_2_c12 <= tile_23_filtered_output_c12(10);
   bh86_w68_2_c12 <= tile_23_filtered_output_c12(11);
   bh86_w69_2_c12 <= tile_23_filtered_output_c12(12);
   bh86_w70_2_c12 <= tile_23_filtered_output_c12(13);
   bh86_w71_2_c12 <= tile_23_filtered_output_c12(14);
   bh86_w72_2_c12 <= tile_23_filtered_output_c12(15);
   bh86_w73_2_c12 <= tile_23_filtered_output_c12(16);
   bh86_w74_2_c12 <= tile_23_filtered_output_c12(17);
   bh86_w75_2_c12 <= tile_23_filtered_output_c12(18);
   bh86_w76_2_c12 <= tile_23_filtered_output_c12(19);
   bh86_w77_2_c12 <= tile_23_filtered_output_c12(20);
   bh86_w78_2_c12 <= tile_23_filtered_output_c12(21);
   bh86_w79_2_c12 <= tile_23_filtered_output_c12(22);
   bh86_w80_2_c12 <= tile_23_filtered_output_c12(23);
   bh86_w81_2_c12 <= tile_23_filtered_output_c12(24);
   bh86_w82_2_c12 <= tile_23_filtered_output_c12(25);
   bh86_w83_2_c12 <= tile_23_filtered_output_c12(26);
   bh86_w84_2_c12 <= tile_23_filtered_output_c12(27);
   bh86_w85_2_c12 <= tile_23_filtered_output_c12(28);
   bh86_w86_2_c12 <= tile_23_filtered_output_c12(29);
   bh86_w87_2_c12 <= tile_23_filtered_output_c12(30);
   bh86_w88_2_c12 <= tile_23_filtered_output_c12(31);
   bh86_w89_2_c12 <= tile_23_filtered_output_c12(32);
   bh86_w90_2_c12 <= tile_23_filtered_output_c12(33);
   bh86_w91_1_c12 <= tile_23_filtered_output_c12(34);
   bh86_w92_1_c12 <= tile_23_filtered_output_c12(35);
   bh86_w93_1_c12 <= tile_23_filtered_output_c12(36);
   bh86_w94_1_c12 <= tile_23_filtered_output_c12(37);
   bh86_w95_1_c12 <= tile_23_filtered_output_c12(38);
   bh86_w96_1_c12 <= tile_23_filtered_output_c12(39);
   bh86_w97_1_c12 <= tile_23_filtered_output_c12(40);
   tile_24_X_c11 <= X(32 downto 16);
   tile_24_Y_c0 <= Y(47 downto 24);
   tile_24_mult: DSPBlock_17x24_Freq300_uid172
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 X => tile_24_X_c11,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c12);

   tile_24_filtered_output_c12 <= unsigned(tile_24_output_c12(40 downto 0));
   bh86_w40_1_c12 <= tile_24_filtered_output_c12(0);
   bh86_w41_1_c12 <= tile_24_filtered_output_c12(1);
   bh86_w42_1_c12 <= tile_24_filtered_output_c12(2);
   bh86_w43_1_c12 <= tile_24_filtered_output_c12(3);
   bh86_w44_13_c12 <= tile_24_filtered_output_c12(4);
   bh86_w45_8_c12 <= tile_24_filtered_output_c12(5);
   bh86_w46_8_c12 <= tile_24_filtered_output_c12(6);
   bh86_w47_9_c12 <= tile_24_filtered_output_c12(7);
   bh86_w48_8_c12 <= tile_24_filtered_output_c12(8);
   bh86_w49_7_c12 <= tile_24_filtered_output_c12(9);
   bh86_w50_8_c12 <= tile_24_filtered_output_c12(10);
   bh86_w51_6_c12 <= tile_24_filtered_output_c12(11);
   bh86_w52_6_c12 <= tile_24_filtered_output_c12(12);
   bh86_w53_5_c12 <= tile_24_filtered_output_c12(13);
   bh86_w54_4_c12 <= tile_24_filtered_output_c12(14);
   bh86_w55_3_c12 <= tile_24_filtered_output_c12(15);
   bh86_w56_3_c12 <= tile_24_filtered_output_c12(16);
   bh86_w57_3_c12 <= tile_24_filtered_output_c12(17);
   bh86_w58_3_c12 <= tile_24_filtered_output_c12(18);
   bh86_w59_3_c12 <= tile_24_filtered_output_c12(19);
   bh86_w60_3_c12 <= tile_24_filtered_output_c12(20);
   bh86_w61_3_c12 <= tile_24_filtered_output_c12(21);
   bh86_w62_3_c12 <= tile_24_filtered_output_c12(22);
   bh86_w63_3_c12 <= tile_24_filtered_output_c12(23);
   bh86_w64_3_c12 <= tile_24_filtered_output_c12(24);
   bh86_w65_3_c12 <= tile_24_filtered_output_c12(25);
   bh86_w66_3_c12 <= tile_24_filtered_output_c12(26);
   bh86_w67_3_c12 <= tile_24_filtered_output_c12(27);
   bh86_w68_3_c12 <= tile_24_filtered_output_c12(28);
   bh86_w69_3_c12 <= tile_24_filtered_output_c12(29);
   bh86_w70_3_c12 <= tile_24_filtered_output_c12(30);
   bh86_w71_3_c12 <= tile_24_filtered_output_c12(31);
   bh86_w72_3_c12 <= tile_24_filtered_output_c12(32);
   bh86_w73_3_c12 <= tile_24_filtered_output_c12(33);
   bh86_w74_3_c12 <= tile_24_filtered_output_c12(34);
   bh86_w75_3_c12 <= tile_24_filtered_output_c12(35);
   bh86_w76_3_c12 <= tile_24_filtered_output_c12(36);
   bh86_w77_3_c12 <= tile_24_filtered_output_c12(37);
   bh86_w78_3_c12 <= tile_24_filtered_output_c12(38);
   bh86_w79_3_c12 <= tile_24_filtered_output_c12(39);
   bh86_w80_3_c12 <= tile_24_filtered_output_c12(40);
   tile_25_X_c11 <= X(15 downto 15);
   tile_25_Y_c0 <= Y(29 downto 29);
   tile_25_mult: IntMultiplierLUT_1x1_Freq300_uid174
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_25_X_c11,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c11);

   tile_25_filtered_output_c11 <= unsigned(tile_25_output_c11(0 downto 0));
   bh86_w44_14_c11 <= tile_25_filtered_output_c11(0);
   tile_26_X_c11 <= X(13 downto 13);
   tile_26_Y_c0 <= Y(31 downto 31);
   tile_26_mult: IntMultiplierLUT_1x1_Freq300_uid176
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_26_X_c11,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c11);

   tile_26_filtered_output_c11 <= unsigned(tile_26_output_c11(0 downto 0));
   bh86_w44_15_c11 <= tile_26_filtered_output_c11(0);
   tile_27_X_c11 <= X(15 downto 14);
   tile_27_Y_c0 <= Y(31 downto 30);
   tile_27_mult: IntMultiplierLUT_2x2_Freq300_uid178
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_27_X_c11,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c11);

   tile_27_filtered_output_c11 <= unsigned(tile_27_output_c11(3 downto 0));
   bh86_w44_16_c11 <= tile_27_filtered_output_c11(0);
   bh86_w45_9_c11 <= tile_27_filtered_output_c11(1);
   bh86_w46_9_c11 <= tile_27_filtered_output_c11(2);
   bh86_w47_10_c11 <= tile_27_filtered_output_c11(3);
   tile_28_X_c11 <= X(12 downto 12);
   tile_28_Y_c0 <= Y(32 downto 32);
   tile_28_mult: IntMultiplierLUT_1x1_Freq300_uid183
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_28_X_c11,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c11);

   tile_28_filtered_output_c11 <= unsigned(tile_28_output_c11(0 downto 0));
   bh86_w44_17_c11 <= tile_28_filtered_output_c11(0);
   tile_29_X_c11 <= X(12 downto 11);
   tile_29_Y_c0 <= Y(33 downto 33);
   tile_29_mult: IntMultiplierLUT_2x1_Freq300_uid185
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_29_X_c11,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c11);

   tile_29_filtered_output_c11 <= unsigned(tile_29_output_c11(1 downto 0));
   bh86_w44_18_c11 <= tile_29_filtered_output_c11(0);
   bh86_w45_10_c11 <= tile_29_filtered_output_c11(1);
   tile_30_X_c11 <= X(15 downto 13);
   tile_30_Y_c0 <= Y(33 downto 32);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid187
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_30_X_c11,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c11);

   tile_30_filtered_output_c11 <= unsigned(tile_30_output_c11(4 downto 0));
   bh86_w45_11_c11 <= tile_30_filtered_output_c11(0);
   bh86_w46_10_c11 <= tile_30_filtered_output_c11(1);
   bh86_w47_11_c11 <= tile_30_filtered_output_c11(2);
   bh86_w48_9_c11 <= tile_30_filtered_output_c11(3);
   bh86_w49_8_c11 <= tile_30_filtered_output_c11(4);
   tile_31_X_c11 <= X(9 downto 9);
   tile_31_Y_c0 <= Y(35 downto 35);
   tile_31_mult: IntMultiplierLUT_1x1_Freq300_uid192
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_31_X_c11,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c11);

   tile_31_filtered_output_c11 <= unsigned(tile_31_output_c11(0 downto 0));
   bh86_w44_19_c11 <= tile_31_filtered_output_c11(0);
   tile_32_X_c11 <= X(12 downto 10);
   tile_32_Y_c0 <= Y(35 downto 34);
   tile_32_mult: IntMultiplierLUT_3x2_Freq300_uid194
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_32_X_c11,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c11);

   tile_32_filtered_output_c11 <= unsigned(tile_32_output_c11(4 downto 0));
   bh86_w44_20_c11 <= tile_32_filtered_output_c11(0);
   bh86_w45_12_c11 <= tile_32_filtered_output_c11(1);
   bh86_w46_11_c11 <= tile_32_filtered_output_c11(2);
   bh86_w47_12_c11 <= tile_32_filtered_output_c11(3);
   bh86_w48_10_c11 <= tile_32_filtered_output_c11(4);
   tile_33_X_c11 <= X(15 downto 13);
   tile_33_Y_c0 <= Y(35 downto 34);
   tile_33_mult: IntMultiplierLUT_3x2_Freq300_uid199
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_33_X_c11,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c11);

   tile_33_filtered_output_c11 <= unsigned(tile_33_output_c11(4 downto 0));
   bh86_w47_13_c11 <= tile_33_filtered_output_c11(0);
   bh86_w48_11_c11 <= tile_33_filtered_output_c11(1);
   bh86_w49_9_c11 <= tile_33_filtered_output_c11(2);
   bh86_w50_9_c11 <= tile_33_filtered_output_c11(3);
   bh86_w51_7_c11 <= tile_33_filtered_output_c11(4);
   tile_34_X_c11 <= X(7 downto 7);
   tile_34_Y_c0 <= Y(37 downto 37);
   tile_34_mult: IntMultiplierLUT_1x1_Freq300_uid204
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_34_X_c11,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c11);

   tile_34_filtered_output_c11 <= unsigned(tile_34_output_c11(0 downto 0));
   bh86_w44_21_c11 <= tile_34_filtered_output_c11(0);
   tile_35_X_c11 <= X(9 downto 8);
   tile_35_Y_c0 <= Y(37 downto 36);
   tile_35_mult: IntMultiplierLUT_2x2_Freq300_uid206
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_35_X_c11,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c11);

   tile_35_filtered_output_c11 <= unsigned(tile_35_output_c11(3 downto 0));
   bh86_w44_22_c11 <= tile_35_filtered_output_c11(0);
   bh86_w45_13_c11 <= tile_35_filtered_output_c11(1);
   bh86_w46_12_c11 <= tile_35_filtered_output_c11(2);
   bh86_w47_14_c11 <= tile_35_filtered_output_c11(3);
   tile_36_X_c11 <= X(12 downto 10);
   tile_36_Y_c0 <= Y(37 downto 36);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid211
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_36_X_c11,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c11);

   tile_36_filtered_output_c11 <= unsigned(tile_36_output_c11(4 downto 0));
   bh86_w46_13_c11 <= tile_36_filtered_output_c11(0);
   bh86_w47_15_c11 <= tile_36_filtered_output_c11(1);
   bh86_w48_12_c11 <= tile_36_filtered_output_c11(2);
   bh86_w49_10_c11 <= tile_36_filtered_output_c11(3);
   bh86_w50_10_c11 <= tile_36_filtered_output_c11(4);
   tile_37_X_c11 <= X(15 downto 13);
   tile_37_Y_c0 <= Y(37 downto 36);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid216
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_37_X_c11,
                 Y => tile_37_Y_c0,
                 R => tile_37_output_c11);

   tile_37_filtered_output_c11 <= unsigned(tile_37_output_c11(4 downto 0));
   bh86_w49_11_c11 <= tile_37_filtered_output_c11(0);
   bh86_w50_11_c11 <= tile_37_filtered_output_c11(1);
   bh86_w51_8_c11 <= tile_37_filtered_output_c11(2);
   bh86_w52_7_c11 <= tile_37_filtered_output_c11(3);
   bh86_w53_6_c11 <= tile_37_filtered_output_c11(4);
   tile_38_X_c11 <= X(6 downto 6);
   tile_38_Y_c0 <= Y(38 downto 38);
   tile_38_mult: IntMultiplierLUT_1x1_Freq300_uid221
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_38_X_c11,
                 Y => tile_38_Y_c0,
                 R => tile_38_output_c11);

   tile_38_filtered_output_c11 <= unsigned(tile_38_output_c11(0 downto 0));
   bh86_w44_23_c11 <= tile_38_filtered_output_c11(0);
   tile_39_X_c11 <= X(6 downto 5);
   tile_39_Y_c0 <= Y(39 downto 39);
   tile_39_mult: IntMultiplierLUT_2x1_Freq300_uid223
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_39_X_c11,
                 Y => tile_39_Y_c0,
                 R => tile_39_output_c11);

   tile_39_filtered_output_c11 <= unsigned(tile_39_output_c11(1 downto 0));
   bh86_w44_24_c11 <= tile_39_filtered_output_c11(0);
   bh86_w45_14_c11 <= tile_39_filtered_output_c11(1);
   tile_40_X_c11 <= X(9 downto 7);
   tile_40_Y_c0 <= Y(39 downto 38);
   tile_40_mult: IntMultiplierLUT_3x2_Freq300_uid225
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_40_X_c11,
                 Y => tile_40_Y_c0,
                 R => tile_40_output_c11);

   tile_40_filtered_output_c11 <= unsigned(tile_40_output_c11(4 downto 0));
   bh86_w45_15_c11 <= tile_40_filtered_output_c11(0);
   bh86_w46_14_c11 <= tile_40_filtered_output_c11(1);
   bh86_w47_16_c11 <= tile_40_filtered_output_c11(2);
   bh86_w48_13_c11 <= tile_40_filtered_output_c11(3);
   bh86_w49_12_c11 <= tile_40_filtered_output_c11(4);
   tile_41_X_c11 <= X(12 downto 10);
   tile_41_Y_c0 <= Y(39 downto 38);
   tile_41_mult: IntMultiplierLUT_3x2_Freq300_uid230
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_41_X_c11,
                 Y => tile_41_Y_c0,
                 R => tile_41_output_c11);

   tile_41_filtered_output_c11 <= unsigned(tile_41_output_c11(4 downto 0));
   bh86_w48_14_c11 <= tile_41_filtered_output_c11(0);
   bh86_w49_13_c11 <= tile_41_filtered_output_c11(1);
   bh86_w50_12_c11 <= tile_41_filtered_output_c11(2);
   bh86_w51_9_c11 <= tile_41_filtered_output_c11(3);
   bh86_w52_8_c11 <= tile_41_filtered_output_c11(4);
   tile_42_X_c11 <= X(15 downto 13);
   tile_42_Y_c0 <= Y(39 downto 38);
   tile_42_mult: IntMultiplierLUT_3x2_Freq300_uid235
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_42_X_c11,
                 Y => tile_42_Y_c0,
                 R => tile_42_output_c11);

   tile_42_filtered_output_c11 <= unsigned(tile_42_output_c11(4 downto 0));
   bh86_w51_10_c11 <= tile_42_filtered_output_c11(0);
   bh86_w52_9_c11 <= tile_42_filtered_output_c11(1);
   bh86_w53_7_c11 <= tile_42_filtered_output_c11(2);
   bh86_w54_5_c11 <= tile_42_filtered_output_c11(3);
   bh86_w55_4_c11 <= tile_42_filtered_output_c11(4);
   tile_43_X_c11 <= X(3 downto 3);
   tile_43_Y_c0 <= Y(41 downto 41);
   tile_43_mult: IntMultiplierLUT_1x1_Freq300_uid240
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_43_X_c11,
                 Y => tile_43_Y_c0,
                 R => tile_43_output_c11);

   tile_43_filtered_output_c11 <= unsigned(tile_43_output_c11(0 downto 0));
   bh86_w44_25_c11 <= tile_43_filtered_output_c11(0);
   tile_44_X_c11 <= X(6 downto 4);
   tile_44_Y_c0 <= Y(41 downto 40);
   tile_44_mult: IntMultiplierLUT_3x2_Freq300_uid242
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_44_X_c11,
                 Y => tile_44_Y_c0,
                 R => tile_44_output_c11);

   tile_44_filtered_output_c11 <= unsigned(tile_44_output_c11(4 downto 0));
   bh86_w44_26_c11 <= tile_44_filtered_output_c11(0);
   bh86_w45_16_c11 <= tile_44_filtered_output_c11(1);
   bh86_w46_15_c11 <= tile_44_filtered_output_c11(2);
   bh86_w47_17_c11 <= tile_44_filtered_output_c11(3);
   bh86_w48_15_c11 <= tile_44_filtered_output_c11(4);
   tile_45_X_c11 <= X(9 downto 7);
   tile_45_Y_c0 <= Y(41 downto 40);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid247
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_45_X_c11,
                 Y => tile_45_Y_c0,
                 R => tile_45_output_c11);

   tile_45_filtered_output_c11 <= unsigned(tile_45_output_c11(4 downto 0));
   bh86_w47_18_c11 <= tile_45_filtered_output_c11(0);
   bh86_w48_16_c11 <= tile_45_filtered_output_c11(1);
   bh86_w49_14_c11 <= tile_45_filtered_output_c11(2);
   bh86_w50_13_c11 <= tile_45_filtered_output_c11(3);
   bh86_w51_11_c11 <= tile_45_filtered_output_c11(4);
   tile_46_X_c11 <= X(12 downto 10);
   tile_46_Y_c0 <= Y(41 downto 40);
   tile_46_mult: IntMultiplierLUT_3x2_Freq300_uid252
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_46_X_c11,
                 Y => tile_46_Y_c0,
                 R => tile_46_output_c11);

   tile_46_filtered_output_c11 <= unsigned(tile_46_output_c11(4 downto 0));
   bh86_w50_14_c11 <= tile_46_filtered_output_c11(0);
   bh86_w51_12_c11 <= tile_46_filtered_output_c11(1);
   bh86_w52_10_c11 <= tile_46_filtered_output_c11(2);
   bh86_w53_8_c11 <= tile_46_filtered_output_c11(3);
   bh86_w54_6_c11 <= tile_46_filtered_output_c11(4);
   tile_47_X_c11 <= X(15 downto 13);
   tile_47_Y_c0 <= Y(41 downto 40);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid257
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_47_X_c11,
                 Y => tile_47_Y_c0,
                 R => tile_47_output_c11);

   tile_47_filtered_output_c11 <= unsigned(tile_47_output_c11(4 downto 0));
   bh86_w53_9_c11 <= tile_47_filtered_output_c11(0);
   bh86_w54_7_c11 <= tile_47_filtered_output_c11(1);
   bh86_w55_5_c11 <= tile_47_filtered_output_c11(2);
   bh86_w56_4_c11 <= tile_47_filtered_output_c11(3);
   bh86_w57_4_c11 <= tile_47_filtered_output_c11(4);
   tile_48_X_c11 <= X(1 downto 1);
   tile_48_Y_c0 <= Y(43 downto 43);
   tile_48_mult: IntMultiplierLUT_1x1_Freq300_uid262
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_48_X_c11,
                 Y => tile_48_Y_c0,
                 R => tile_48_output_c11);

   tile_48_filtered_output_c11 <= unsigned(tile_48_output_c11(0 downto 0));
   bh86_w44_27_c11 <= tile_48_filtered_output_c11(0);
   tile_49_X_c11 <= X(3 downto 2);
   tile_49_Y_c0 <= Y(43 downto 42);
   tile_49_mult: IntMultiplierLUT_2x2_Freq300_uid264
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_49_X_c11,
                 Y => tile_49_Y_c0,
                 R => tile_49_output_c11);

   tile_49_filtered_output_c11 <= unsigned(tile_49_output_c11(3 downto 0));
   bh86_w44_28_c11 <= tile_49_filtered_output_c11(0);
   bh86_w45_17_c11 <= tile_49_filtered_output_c11(1);
   bh86_w46_16_c11 <= tile_49_filtered_output_c11(2);
   bh86_w47_19_c11 <= tile_49_filtered_output_c11(3);
   tile_50_X_c11 <= X(6 downto 4);
   tile_50_Y_c0 <= Y(43 downto 42);
   tile_50_mult: IntMultiplierLUT_3x2_Freq300_uid269
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_50_X_c11,
                 Y => tile_50_Y_c0,
                 R => tile_50_output_c11);

   tile_50_filtered_output_c11 <= unsigned(tile_50_output_c11(4 downto 0));
   bh86_w46_17_c11 <= tile_50_filtered_output_c11(0);
   bh86_w47_20_c11 <= tile_50_filtered_output_c11(1);
   bh86_w48_17_c11 <= tile_50_filtered_output_c11(2);
   bh86_w49_15_c11 <= tile_50_filtered_output_c11(3);
   bh86_w50_15_c11 <= tile_50_filtered_output_c11(4);
   tile_51_X_c11 <= X(9 downto 7);
   tile_51_Y_c0 <= Y(43 downto 42);
   tile_51_mult: IntMultiplierLUT_3x2_Freq300_uid274
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_51_X_c11,
                 Y => tile_51_Y_c0,
                 R => tile_51_output_c11);

   tile_51_filtered_output_c11 <= unsigned(tile_51_output_c11(4 downto 0));
   bh86_w49_16_c11 <= tile_51_filtered_output_c11(0);
   bh86_w50_16_c11 <= tile_51_filtered_output_c11(1);
   bh86_w51_13_c11 <= tile_51_filtered_output_c11(2);
   bh86_w52_11_c11 <= tile_51_filtered_output_c11(3);
   bh86_w53_10_c11 <= tile_51_filtered_output_c11(4);
   tile_52_X_c11 <= X(12 downto 10);
   tile_52_Y_c0 <= Y(43 downto 42);
   tile_52_mult: IntMultiplierLUT_3x2_Freq300_uid279
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_52_X_c11,
                 Y => tile_52_Y_c0,
                 R => tile_52_output_c11);

   tile_52_filtered_output_c11 <= unsigned(tile_52_output_c11(4 downto 0));
   bh86_w52_12_c11 <= tile_52_filtered_output_c11(0);
   bh86_w53_11_c11 <= tile_52_filtered_output_c11(1);
   bh86_w54_8_c11 <= tile_52_filtered_output_c11(2);
   bh86_w55_6_c11 <= tile_52_filtered_output_c11(3);
   bh86_w56_5_c11 <= tile_52_filtered_output_c11(4);
   tile_53_X_c11 <= X(15 downto 13);
   tile_53_Y_c0 <= Y(43 downto 42);
   tile_53_mult: IntMultiplierLUT_3x2_Freq300_uid284
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_53_X_c11,
                 Y => tile_53_Y_c0,
                 R => tile_53_output_c11);

   tile_53_filtered_output_c11 <= unsigned(tile_53_output_c11(4 downto 0));
   bh86_w55_7_c11 <= tile_53_filtered_output_c11(0);
   bh86_w56_6_c11 <= tile_53_filtered_output_c11(1);
   bh86_w57_5_c11 <= tile_53_filtered_output_c11(2);
   bh86_w58_4_c11 <= tile_53_filtered_output_c11(3);
   bh86_w59_4_c11 <= tile_53_filtered_output_c11(4);
   tile_54_X_c11 <= X(0 downto 0);
   tile_54_Y_c0 <= Y(45 downto 44);
   tile_54_mult: IntMultiplierLUT_1x2_Freq300_uid289
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_54_X_c11,
                 Y => tile_54_Y_c0,
                 R => tile_54_output_c11);

   tile_54_filtered_output_c11 <= unsigned(tile_54_output_c11(1 downto 0));
   bh86_w44_29_c11 <= tile_54_filtered_output_c11(0);
   bh86_w45_18_c11 <= tile_54_filtered_output_c11(1);
   tile_55_X_c11 <= X(3 downto 1);
   tile_55_Y_c0 <= Y(45 downto 44);
   tile_55_mult: IntMultiplierLUT_3x2_Freq300_uid291
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_55_X_c11,
                 Y => tile_55_Y_c0,
                 R => tile_55_output_c11);

   tile_55_filtered_output_c11 <= unsigned(tile_55_output_c11(4 downto 0));
   bh86_w45_19_c11 <= tile_55_filtered_output_c11(0);
   bh86_w46_18_c11 <= tile_55_filtered_output_c11(1);
   bh86_w47_21_c11 <= tile_55_filtered_output_c11(2);
   bh86_w48_18_c11 <= tile_55_filtered_output_c11(3);
   bh86_w49_17_c11 <= tile_55_filtered_output_c11(4);
   tile_56_X_c11 <= X(6 downto 4);
   tile_56_Y_c0 <= Y(45 downto 44);
   tile_56_mult: IntMultiplierLUT_3x2_Freq300_uid296
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_56_X_c11,
                 Y => tile_56_Y_c0,
                 R => tile_56_output_c11);

   tile_56_filtered_output_c11 <= unsigned(tile_56_output_c11(4 downto 0));
   bh86_w48_19_c11 <= tile_56_filtered_output_c11(0);
   bh86_w49_18_c11 <= tile_56_filtered_output_c11(1);
   bh86_w50_17_c11 <= tile_56_filtered_output_c11(2);
   bh86_w51_14_c11 <= tile_56_filtered_output_c11(3);
   bh86_w52_13_c11 <= tile_56_filtered_output_c11(4);
   tile_57_X_c11 <= X(9 downto 7);
   tile_57_Y_c0 <= Y(45 downto 44);
   tile_57_mult: IntMultiplierLUT_3x2_Freq300_uid301
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_57_X_c11,
                 Y => tile_57_Y_c0,
                 R => tile_57_output_c11);

   tile_57_filtered_output_c11 <= unsigned(tile_57_output_c11(4 downto 0));
   bh86_w51_15_c11 <= tile_57_filtered_output_c11(0);
   bh86_w52_14_c11 <= tile_57_filtered_output_c11(1);
   bh86_w53_12_c11 <= tile_57_filtered_output_c11(2);
   bh86_w54_9_c11 <= tile_57_filtered_output_c11(3);
   bh86_w55_8_c11 <= tile_57_filtered_output_c11(4);
   tile_58_X_c11 <= X(12 downto 10);
   tile_58_Y_c0 <= Y(45 downto 44);
   tile_58_mult: IntMultiplierLUT_3x2_Freq300_uid306
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_58_X_c11,
                 Y => tile_58_Y_c0,
                 R => tile_58_output_c11);

   tile_58_filtered_output_c11 <= unsigned(tile_58_output_c11(4 downto 0));
   bh86_w54_10_c11 <= tile_58_filtered_output_c11(0);
   bh86_w55_9_c11 <= tile_58_filtered_output_c11(1);
   bh86_w56_7_c11 <= tile_58_filtered_output_c11(2);
   bh86_w57_6_c11 <= tile_58_filtered_output_c11(3);
   bh86_w58_5_c11 <= tile_58_filtered_output_c11(4);
   tile_59_X_c11 <= X(15 downto 13);
   tile_59_Y_c0 <= Y(45 downto 44);
   tile_59_mult: IntMultiplierLUT_3x2_Freq300_uid311
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_59_X_c11,
                 Y => tile_59_Y_c0,
                 R => tile_59_output_c11);

   tile_59_filtered_output_c11 <= unsigned(tile_59_output_c11(4 downto 0));
   bh86_w57_7_c11 <= tile_59_filtered_output_c11(0);
   bh86_w58_6_c11 <= tile_59_filtered_output_c11(1);
   bh86_w59_5_c11 <= tile_59_filtered_output_c11(2);
   bh86_w60_4_c11 <= tile_59_filtered_output_c11(3);
   bh86_w61_4_c11 <= tile_59_filtered_output_c11(4);
   tile_60_X_c11 <= X(0 downto 0);
   tile_60_Y_c0 <= Y(47 downto 46);
   tile_60_mult: IntMultiplierLUT_1x2_Freq300_uid316
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_60_X_c11,
                 Y => tile_60_Y_c0,
                 R => tile_60_output_c11);

   tile_60_filtered_output_c11 <= unsigned(tile_60_output_c11(1 downto 0));
   bh86_w46_19_c11 <= tile_60_filtered_output_c11(0);
   bh86_w47_22_c11 <= tile_60_filtered_output_c11(1);
   tile_61_X_c11 <= X(3 downto 1);
   tile_61_Y_c0 <= Y(47 downto 46);
   tile_61_mult: IntMultiplierLUT_3x2_Freq300_uid318
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_61_X_c11,
                 Y => tile_61_Y_c0,
                 R => tile_61_output_c11);

   tile_61_filtered_output_c11 <= unsigned(tile_61_output_c11(4 downto 0));
   bh86_w47_23_c11 <= tile_61_filtered_output_c11(0);
   bh86_w48_20_c11 <= tile_61_filtered_output_c11(1);
   bh86_w49_19_c11 <= tile_61_filtered_output_c11(2);
   bh86_w50_18_c11 <= tile_61_filtered_output_c11(3);
   bh86_w51_16_c11 <= tile_61_filtered_output_c11(4);
   tile_62_X_c11 <= X(6 downto 4);
   tile_62_Y_c0 <= Y(47 downto 46);
   tile_62_mult: IntMultiplierLUT_3x2_Freq300_uid323
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_62_X_c11,
                 Y => tile_62_Y_c0,
                 R => tile_62_output_c11);

   tile_62_filtered_output_c11 <= unsigned(tile_62_output_c11(4 downto 0));
   bh86_w50_19_c11 <= tile_62_filtered_output_c11(0);
   bh86_w51_17_c11 <= tile_62_filtered_output_c11(1);
   bh86_w52_15_c11 <= tile_62_filtered_output_c11(2);
   bh86_w53_13_c11 <= tile_62_filtered_output_c11(3);
   bh86_w54_11_c11 <= tile_62_filtered_output_c11(4);
   tile_63_X_c11 <= X(9 downto 7);
   tile_63_Y_c0 <= Y(47 downto 46);
   tile_63_mult: IntMultiplierLUT_3x2_Freq300_uid328
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_63_X_c11,
                 Y => tile_63_Y_c0,
                 R => tile_63_output_c11);

   tile_63_filtered_output_c11 <= unsigned(tile_63_output_c11(4 downto 0));
   bh86_w53_14_c11 <= tile_63_filtered_output_c11(0);
   bh86_w54_12_c11 <= tile_63_filtered_output_c11(1);
   bh86_w55_10_c11 <= tile_63_filtered_output_c11(2);
   bh86_w56_8_c11 <= tile_63_filtered_output_c11(3);
   bh86_w57_8_c11 <= tile_63_filtered_output_c11(4);
   tile_64_X_c11 <= X(12 downto 10);
   tile_64_Y_c0 <= Y(47 downto 46);
   tile_64_mult: IntMultiplierLUT_3x2_Freq300_uid333
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_64_X_c11,
                 Y => tile_64_Y_c0,
                 R => tile_64_output_c11);

   tile_64_filtered_output_c11 <= unsigned(tile_64_output_c11(4 downto 0));
   bh86_w56_9_c11 <= tile_64_filtered_output_c11(0);
   bh86_w57_9_c11 <= tile_64_filtered_output_c11(1);
   bh86_w58_7_c11 <= tile_64_filtered_output_c11(2);
   bh86_w59_6_c11 <= tile_64_filtered_output_c11(3);
   bh86_w60_5_c11 <= tile_64_filtered_output_c11(4);
   tile_65_X_c11 <= X(15 downto 13);
   tile_65_Y_c0 <= Y(47 downto 46);
   tile_65_mult: IntMultiplierLUT_3x2_Freq300_uid338
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_65_X_c11,
                 Y => tile_65_Y_c0,
                 R => tile_65_output_c11);

   tile_65_filtered_output_c11 <= unsigned(tile_65_output_c11(4 downto 0));
   bh86_w59_7_c11 <= tile_65_filtered_output_c11(0);
   bh86_w60_6_c11 <= tile_65_filtered_output_c11(1);
   bh86_w61_5_c11 <= tile_65_filtered_output_c11(2);
   bh86_w62_4_c11 <= tile_65_filtered_output_c11(3);
   bh86_w63_4_c11 <= tile_65_filtered_output_c11(4);
   tile_66_X_c11 <= X(50 downto 50);
   tile_66_Y_c0 <= Y(48 downto 48);
   tile_66_mult: IntMultiplierLUT_1x1_Freq300_uid343
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_66_X_c11,
                 Y => tile_66_Y_c0,
                 R => tile_66_output_c11);

   tile_66_filtered_output_c11 <= unsigned(tile_66_output_c11(0 downto 0));
   bh86_w98_1_c11 <= tile_66_filtered_output_c11(0);
   tile_67_X_c11 <= X(54 downto 51);
   tile_67_Y_c0 <= Y(48 downto 48);
   tile_67_mult: IntMultiplierLUT_4x1_Freq300_uid345
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_67_X_c11,
                 Y => tile_67_Y_c0,
                 R => tile_67_output_c11);

   tile_67_filtered_output_c11 <= unsigned(tile_67_output_c11(3 downto 0));
   bh86_w99_1_c11 <= tile_67_filtered_output_c11(0);
   bh86_w100_1_c11 <= tile_67_filtered_output_c11(1);
   bh86_w101_1_c11 <= tile_67_filtered_output_c11(2);
   bh86_w102_1_c11 <= tile_67_filtered_output_c11(3);
   tile_68_X_c11 <= X(58 downto 55);
   tile_68_Y_c0 <= Y(48 downto 48);
   tile_68_mult: IntMultiplierLUT_4x1_Freq300_uid347
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_68_X_c11,
                 Y => tile_68_Y_c0,
                 R => tile_68_output_c11);

   tile_68_filtered_output_c11 <= unsigned(tile_68_output_c11(3 downto 0));
   bh86_w103_1_c11 <= tile_68_filtered_output_c11(0);
   bh86_w104_1_c11 <= tile_68_filtered_output_c11(1);
   bh86_w105_1_c11 <= tile_68_filtered_output_c11(2);
   bh86_w106_1_c11 <= tile_68_filtered_output_c11(3);
   tile_69_X_c11 <= X(62 downto 59);
   tile_69_Y_c0 <= Y(48 downto 48);
   tile_69_mult: IntMultiplierLUT_4x1_Freq300_uid349
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_69_X_c11,
                 Y => tile_69_Y_c0,
                 R => tile_69_output_c11);

   tile_69_filtered_output_c11 <= unsigned(tile_69_output_c11(3 downto 0));
   bh86_w107_1_c11 <= tile_69_filtered_output_c11(0);
   bh86_w108_1_c11 <= tile_69_filtered_output_c11(1);
   bh86_w109_1_c11 <= tile_69_filtered_output_c11(2);
   bh86_w110_1_c11 <= tile_69_filtered_output_c11(3);
   tile_70_X_c11 <= X(66 downto 63);
   tile_70_Y_c0 <= Y(48 downto 48);
   tile_70_mult: IntMultiplierLUT_4x1_Freq300_uid351
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_70_X_c11,
                 Y => tile_70_Y_c0,
                 R => tile_70_output_c11);

   tile_70_filtered_output_c11 <= unsigned(tile_70_output_c11(3 downto 0));
   bh86_w111_1_c11 <= tile_70_filtered_output_c11(0);
   bh86_w112_1_c11 <= tile_70_filtered_output_c11(1);
   bh86_w113_1_c11 <= tile_70_filtered_output_c11(2);
   bh86_w114_1_c11 <= tile_70_filtered_output_c11(3);
   tile_71_X_c11 <= X(51 downto 50);
   tile_71_Y_c0 <= Y(50 downto 49);
   tile_71_mult: IntMultiplierLUT_2x2_Freq300_uid353
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_71_X_c11,
                 Y => tile_71_Y_c0,
                 R => tile_71_output_c11);

   tile_71_filtered_output_c11 <= unsigned(tile_71_output_c11(3 downto 0));
   bh86_w99_2_c11 <= tile_71_filtered_output_c11(0);
   bh86_w100_2_c11 <= tile_71_filtered_output_c11(1);
   bh86_w101_2_c11 <= tile_71_filtered_output_c11(2);
   bh86_w102_2_c11 <= tile_71_filtered_output_c11(3);
   tile_72_X_c11 <= X(54 downto 52);
   tile_72_Y_c0 <= Y(50 downto 49);
   tile_72_mult: IntMultiplierLUT_3x2_Freq300_uid358
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_72_X_c11,
                 Y => tile_72_Y_c0,
                 R => tile_72_output_c11);

   tile_72_filtered_output_c11 <= unsigned(tile_72_output_c11(4 downto 0));
   bh86_w101_3_c11 <= tile_72_filtered_output_c11(0);
   bh86_w102_3_c11 <= tile_72_filtered_output_c11(1);
   bh86_w103_2_c11 <= tile_72_filtered_output_c11(2);
   bh86_w104_2_c11 <= tile_72_filtered_output_c11(3);
   bh86_w105_2_c11 <= tile_72_filtered_output_c11(4);
   tile_73_X_c11 <= X(57 downto 55);
   tile_73_Y_c0 <= Y(50 downto 49);
   tile_73_mult: IntMultiplierLUT_3x2_Freq300_uid363
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_73_X_c11,
                 Y => tile_73_Y_c0,
                 R => tile_73_output_c11);

   tile_73_filtered_output_c11 <= unsigned(tile_73_output_c11(4 downto 0));
   bh86_w104_3_c11 <= tile_73_filtered_output_c11(0);
   bh86_w105_3_c11 <= tile_73_filtered_output_c11(1);
   bh86_w106_2_c11 <= tile_73_filtered_output_c11(2);
   bh86_w107_2_c11 <= tile_73_filtered_output_c11(3);
   bh86_w108_2_c11 <= tile_73_filtered_output_c11(4);
   tile_74_X_c11 <= X(60 downto 58);
   tile_74_Y_c0 <= Y(50 downto 49);
   tile_74_mult: IntMultiplierLUT_3x2_Freq300_uid368
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_74_X_c11,
                 Y => tile_74_Y_c0,
                 R => tile_74_output_c11);

   tile_74_filtered_output_c11 <= unsigned(tile_74_output_c11(4 downto 0));
   bh86_w107_3_c11 <= tile_74_filtered_output_c11(0);
   bh86_w108_3_c11 <= tile_74_filtered_output_c11(1);
   bh86_w109_2_c11 <= tile_74_filtered_output_c11(2);
   bh86_w110_2_c11 <= tile_74_filtered_output_c11(3);
   bh86_w111_2_c11 <= tile_74_filtered_output_c11(4);
   tile_75_X_c11 <= X(63 downto 61);
   tile_75_Y_c0 <= Y(50 downto 49);
   tile_75_mult: IntMultiplierLUT_3x2_Freq300_uid373
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_75_X_c11,
                 Y => tile_75_Y_c0,
                 R => tile_75_output_c11);

   tile_75_filtered_output_c11 <= unsigned(tile_75_output_c11(4 downto 0));
   bh86_w110_3_c11 <= tile_75_filtered_output_c11(0);
   bh86_w111_3_c11 <= tile_75_filtered_output_c11(1);
   bh86_w112_2_c11 <= tile_75_filtered_output_c11(2);
   bh86_w113_2_c11 <= tile_75_filtered_output_c11(3);
   bh86_w114_2_c11 <= tile_75_filtered_output_c11(4);
   tile_76_X_c11 <= X(66 downto 64);
   tile_76_Y_c0 <= Y(50 downto 49);
   tile_76_mult: IntMultiplierLUT_3x2_Freq300_uid378
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_76_X_c11,
                 Y => tile_76_Y_c0,
                 R => tile_76_output_c11);

   tile_76_filtered_output_c11 <= unsigned(tile_76_output_c11(4 downto 0));
   bh86_w113_3_c11 <= tile_76_filtered_output_c11(0);
   bh86_w114_3_c11 <= tile_76_filtered_output_c11(1);
   bh86_w115_0_c11 <= tile_76_filtered_output_c11(2);
   bh86_w116_0_c11 <= tile_76_filtered_output_c11(3);
   bh86_w117_0_c11 <= tile_76_filtered_output_c11(4);
   tile_77_X_c11 <= X(51 downto 50);
   tile_77_Y_c0 <= Y(52 downto 51);
   tile_77_mult: IntMultiplierLUT_2x2_Freq300_uid383
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_77_X_c11,
                 Y => tile_77_Y_c0,
                 R => tile_77_output_c11);

   tile_77_filtered_output_c11 <= unsigned(tile_77_output_c11(3 downto 0));
   bh86_w101_4_c11 <= tile_77_filtered_output_c11(0);
   bh86_w102_4_c11 <= tile_77_filtered_output_c11(1);
   bh86_w103_3_c11 <= tile_77_filtered_output_c11(2);
   bh86_w104_4_c11 <= tile_77_filtered_output_c11(3);
   tile_78_X_c11 <= X(54 downto 52);
   tile_78_Y_c0 <= Y(52 downto 51);
   tile_78_mult: IntMultiplierLUT_3x2_Freq300_uid388
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_78_X_c11,
                 Y => tile_78_Y_c0,
                 R => tile_78_output_c11);

   tile_78_filtered_output_c11 <= unsigned(tile_78_output_c11(4 downto 0));
   bh86_w103_4_c11 <= tile_78_filtered_output_c11(0);
   bh86_w104_5_c11 <= tile_78_filtered_output_c11(1);
   bh86_w105_4_c11 <= tile_78_filtered_output_c11(2);
   bh86_w106_3_c11 <= tile_78_filtered_output_c11(3);
   bh86_w107_4_c11 <= tile_78_filtered_output_c11(4);
   tile_79_X_c11 <= X(57 downto 55);
   tile_79_Y_c0 <= Y(52 downto 51);
   tile_79_mult: IntMultiplierLUT_3x2_Freq300_uid393
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_79_X_c11,
                 Y => tile_79_Y_c0,
                 R => tile_79_output_c11);

   tile_79_filtered_output_c11 <= unsigned(tile_79_output_c11(4 downto 0));
   bh86_w106_4_c11 <= tile_79_filtered_output_c11(0);
   bh86_w107_5_c11 <= tile_79_filtered_output_c11(1);
   bh86_w108_4_c11 <= tile_79_filtered_output_c11(2);
   bh86_w109_3_c11 <= tile_79_filtered_output_c11(3);
   bh86_w110_4_c11 <= tile_79_filtered_output_c11(4);
   tile_80_X_c11 <= X(60 downto 58);
   tile_80_Y_c0 <= Y(52 downto 51);
   tile_80_mult: IntMultiplierLUT_3x2_Freq300_uid398
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_80_X_c11,
                 Y => tile_80_Y_c0,
                 R => tile_80_output_c11);

   tile_80_filtered_output_c11 <= unsigned(tile_80_output_c11(4 downto 0));
   bh86_w109_4_c11 <= tile_80_filtered_output_c11(0);
   bh86_w110_5_c11 <= tile_80_filtered_output_c11(1);
   bh86_w111_4_c11 <= tile_80_filtered_output_c11(2);
   bh86_w112_3_c11 <= tile_80_filtered_output_c11(3);
   bh86_w113_4_c11 <= tile_80_filtered_output_c11(4);
   tile_81_X_c11 <= X(63 downto 61);
   tile_81_Y_c0 <= Y(52 downto 51);
   tile_81_mult: IntMultiplierLUT_3x2_Freq300_uid403
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_81_X_c11,
                 Y => tile_81_Y_c0,
                 R => tile_81_output_c11);

   tile_81_filtered_output_c11 <= unsigned(tile_81_output_c11(4 downto 0));
   bh86_w112_4_c11 <= tile_81_filtered_output_c11(0);
   bh86_w113_5_c11 <= tile_81_filtered_output_c11(1);
   bh86_w114_4_c11 <= tile_81_filtered_output_c11(2);
   bh86_w115_1_c11 <= tile_81_filtered_output_c11(3);
   bh86_w116_1_c11 <= tile_81_filtered_output_c11(4);
   tile_82_X_c11 <= X(66 downto 64);
   tile_82_Y_c0 <= Y(52 downto 51);
   tile_82_mult: IntMultiplierLUT_3x2_Freq300_uid408
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_82_X_c11,
                 Y => tile_82_Y_c0,
                 R => tile_82_output_c11);

   tile_82_filtered_output_c11 <= unsigned(tile_82_output_c11(4 downto 0));
   bh86_w115_2_c11 <= tile_82_filtered_output_c11(0);
   bh86_w116_2_c11 <= tile_82_filtered_output_c11(1);
   bh86_w117_1_c11 <= tile_82_filtered_output_c11(2);
   bh86_w118_0_c11 <= tile_82_filtered_output_c11(3);
   bh86_w119_0_c11 <= tile_82_filtered_output_c11(4);
   tile_83_X_c11 <= X(33 downto 33);
   tile_83_Y_c0 <= Y(48 downto 48);
   tile_83_mult: IntMultiplierLUT_1x1_Freq300_uid413
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_83_X_c11,
                 Y => tile_83_Y_c0,
                 R => tile_83_output_c11);

   tile_83_filtered_output_c11 <= unsigned(tile_83_output_c11(0 downto 0));
   bh86_w81_3_c11 <= tile_83_filtered_output_c11(0);
   tile_84_X_c11 <= X(37 downto 34);
   tile_84_Y_c0 <= Y(48 downto 48);
   tile_84_mult: IntMultiplierLUT_4x1_Freq300_uid415
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_84_X_c11,
                 Y => tile_84_Y_c0,
                 R => tile_84_output_c11);

   tile_84_filtered_output_c11 <= unsigned(tile_84_output_c11(3 downto 0));
   bh86_w82_3_c11 <= tile_84_filtered_output_c11(0);
   bh86_w83_3_c11 <= tile_84_filtered_output_c11(1);
   bh86_w84_3_c11 <= tile_84_filtered_output_c11(2);
   bh86_w85_3_c11 <= tile_84_filtered_output_c11(3);
   tile_85_X_c11 <= X(41 downto 38);
   tile_85_Y_c0 <= Y(48 downto 48);
   tile_85_mult: IntMultiplierLUT_4x1_Freq300_uid417
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_85_X_c11,
                 Y => tile_85_Y_c0,
                 R => tile_85_output_c11);

   tile_85_filtered_output_c11 <= unsigned(tile_85_output_c11(3 downto 0));
   bh86_w86_3_c11 <= tile_85_filtered_output_c11(0);
   bh86_w87_3_c11 <= tile_85_filtered_output_c11(1);
   bh86_w88_3_c11 <= tile_85_filtered_output_c11(2);
   bh86_w89_3_c11 <= tile_85_filtered_output_c11(3);
   tile_86_X_c11 <= X(45 downto 42);
   tile_86_Y_c0 <= Y(48 downto 48);
   tile_86_mult: IntMultiplierLUT_4x1_Freq300_uid419
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_86_X_c11,
                 Y => tile_86_Y_c0,
                 R => tile_86_output_c11);

   tile_86_filtered_output_c11 <= unsigned(tile_86_output_c11(3 downto 0));
   bh86_w90_3_c11 <= tile_86_filtered_output_c11(0);
   bh86_w91_2_c11 <= tile_86_filtered_output_c11(1);
   bh86_w92_2_c11 <= tile_86_filtered_output_c11(2);
   bh86_w93_2_c11 <= tile_86_filtered_output_c11(3);
   tile_87_X_c11 <= X(49 downto 46);
   tile_87_Y_c0 <= Y(48 downto 48);
   tile_87_mult: IntMultiplierLUT_4x1_Freq300_uid421
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_87_X_c11,
                 Y => tile_87_Y_c0,
                 R => tile_87_output_c11);

   tile_87_filtered_output_c11 <= unsigned(tile_87_output_c11(3 downto 0));
   bh86_w94_2_c11 <= tile_87_filtered_output_c11(0);
   bh86_w95_2_c11 <= tile_87_filtered_output_c11(1);
   bh86_w96_2_c11 <= tile_87_filtered_output_c11(2);
   bh86_w97_2_c11 <= tile_87_filtered_output_c11(3);
   tile_88_X_c11 <= X(34 downto 33);
   tile_88_Y_c0 <= Y(50 downto 49);
   tile_88_mult: IntMultiplierLUT_2x2_Freq300_uid423
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_88_X_c11,
                 Y => tile_88_Y_c0,
                 R => tile_88_output_c11);

   tile_88_filtered_output_c11 <= unsigned(tile_88_output_c11(3 downto 0));
   bh86_w82_4_c11 <= tile_88_filtered_output_c11(0);
   bh86_w83_4_c11 <= tile_88_filtered_output_c11(1);
   bh86_w84_4_c11 <= tile_88_filtered_output_c11(2);
   bh86_w85_4_c11 <= tile_88_filtered_output_c11(3);
   tile_89_X_c11 <= X(37 downto 35);
   tile_89_Y_c0 <= Y(50 downto 49);
   tile_89_mult: IntMultiplierLUT_3x2_Freq300_uid428
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_89_X_c11,
                 Y => tile_89_Y_c0,
                 R => tile_89_output_c11);

   tile_89_filtered_output_c11 <= unsigned(tile_89_output_c11(4 downto 0));
   bh86_w84_5_c11 <= tile_89_filtered_output_c11(0);
   bh86_w85_5_c11 <= tile_89_filtered_output_c11(1);
   bh86_w86_4_c11 <= tile_89_filtered_output_c11(2);
   bh86_w87_4_c11 <= tile_89_filtered_output_c11(3);
   bh86_w88_4_c11 <= tile_89_filtered_output_c11(4);
   tile_90_X_c11 <= X(40 downto 38);
   tile_90_Y_c0 <= Y(50 downto 49);
   tile_90_mult: IntMultiplierLUT_3x2_Freq300_uid433
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_90_X_c11,
                 Y => tile_90_Y_c0,
                 R => tile_90_output_c11);

   tile_90_filtered_output_c11 <= unsigned(tile_90_output_c11(4 downto 0));
   bh86_w87_5_c11 <= tile_90_filtered_output_c11(0);
   bh86_w88_5_c11 <= tile_90_filtered_output_c11(1);
   bh86_w89_4_c11 <= tile_90_filtered_output_c11(2);
   bh86_w90_4_c11 <= tile_90_filtered_output_c11(3);
   bh86_w91_3_c11 <= tile_90_filtered_output_c11(4);
   tile_91_X_c11 <= X(43 downto 41);
   tile_91_Y_c0 <= Y(50 downto 49);
   tile_91_mult: IntMultiplierLUT_3x2_Freq300_uid438
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_91_X_c11,
                 Y => tile_91_Y_c0,
                 R => tile_91_output_c11);

   tile_91_filtered_output_c11 <= unsigned(tile_91_output_c11(4 downto 0));
   bh86_w90_5_c11 <= tile_91_filtered_output_c11(0);
   bh86_w91_4_c11 <= tile_91_filtered_output_c11(1);
   bh86_w92_3_c11 <= tile_91_filtered_output_c11(2);
   bh86_w93_3_c11 <= tile_91_filtered_output_c11(3);
   bh86_w94_3_c11 <= tile_91_filtered_output_c11(4);
   tile_92_X_c11 <= X(46 downto 44);
   tile_92_Y_c0 <= Y(50 downto 49);
   tile_92_mult: IntMultiplierLUT_3x2_Freq300_uid443
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_92_X_c11,
                 Y => tile_92_Y_c0,
                 R => tile_92_output_c11);

   tile_92_filtered_output_c11 <= unsigned(tile_92_output_c11(4 downto 0));
   bh86_w93_4_c11 <= tile_92_filtered_output_c11(0);
   bh86_w94_4_c11 <= tile_92_filtered_output_c11(1);
   bh86_w95_3_c11 <= tile_92_filtered_output_c11(2);
   bh86_w96_3_c11 <= tile_92_filtered_output_c11(3);
   bh86_w97_3_c11 <= tile_92_filtered_output_c11(4);
   tile_93_X_c11 <= X(49 downto 47);
   tile_93_Y_c0 <= Y(50 downto 49);
   tile_93_mult: IntMultiplierLUT_3x2_Freq300_uid448
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_93_X_c11,
                 Y => tile_93_Y_c0,
                 R => tile_93_output_c11);

   tile_93_filtered_output_c11 <= unsigned(tile_93_output_c11(4 downto 0));
   bh86_w96_4_c11 <= tile_93_filtered_output_c11(0);
   bh86_w97_4_c11 <= tile_93_filtered_output_c11(1);
   bh86_w98_2_c11 <= tile_93_filtered_output_c11(2);
   bh86_w99_3_c11 <= tile_93_filtered_output_c11(3);
   bh86_w100_3_c11 <= tile_93_filtered_output_c11(4);
   tile_94_X_c11 <= X(34 downto 33);
   tile_94_Y_c0 <= Y(52 downto 51);
   tile_94_mult: IntMultiplierLUT_2x2_Freq300_uid453
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_94_X_c11,
                 Y => tile_94_Y_c0,
                 R => tile_94_output_c11);

   tile_94_filtered_output_c11 <= unsigned(tile_94_output_c11(3 downto 0));
   bh86_w84_6_c11 <= tile_94_filtered_output_c11(0);
   bh86_w85_6_c11 <= tile_94_filtered_output_c11(1);
   bh86_w86_5_c11 <= tile_94_filtered_output_c11(2);
   bh86_w87_6_c11 <= tile_94_filtered_output_c11(3);
   tile_95_X_c11 <= X(37 downto 35);
   tile_95_Y_c0 <= Y(52 downto 51);
   tile_95_mult: IntMultiplierLUT_3x2_Freq300_uid458
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_95_X_c11,
                 Y => tile_95_Y_c0,
                 R => tile_95_output_c11);

   tile_95_filtered_output_c11 <= unsigned(tile_95_output_c11(4 downto 0));
   bh86_w86_6_c11 <= tile_95_filtered_output_c11(0);
   bh86_w87_7_c11 <= tile_95_filtered_output_c11(1);
   bh86_w88_6_c11 <= tile_95_filtered_output_c11(2);
   bh86_w89_5_c11 <= tile_95_filtered_output_c11(3);
   bh86_w90_6_c11 <= tile_95_filtered_output_c11(4);
   tile_96_X_c11 <= X(40 downto 38);
   tile_96_Y_c0 <= Y(52 downto 51);
   tile_96_mult: IntMultiplierLUT_3x2_Freq300_uid463
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_96_X_c11,
                 Y => tile_96_Y_c0,
                 R => tile_96_output_c11);

   tile_96_filtered_output_c11 <= unsigned(tile_96_output_c11(4 downto 0));
   bh86_w89_6_c11 <= tile_96_filtered_output_c11(0);
   bh86_w90_7_c11 <= tile_96_filtered_output_c11(1);
   bh86_w91_5_c11 <= tile_96_filtered_output_c11(2);
   bh86_w92_4_c11 <= tile_96_filtered_output_c11(3);
   bh86_w93_5_c11 <= tile_96_filtered_output_c11(4);
   tile_97_X_c11 <= X(43 downto 41);
   tile_97_Y_c0 <= Y(52 downto 51);
   tile_97_mult: IntMultiplierLUT_3x2_Freq300_uid468
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_97_X_c11,
                 Y => tile_97_Y_c0,
                 R => tile_97_output_c11);

   tile_97_filtered_output_c11 <= unsigned(tile_97_output_c11(4 downto 0));
   bh86_w92_5_c11 <= tile_97_filtered_output_c11(0);
   bh86_w93_6_c11 <= tile_97_filtered_output_c11(1);
   bh86_w94_5_c11 <= tile_97_filtered_output_c11(2);
   bh86_w95_4_c11 <= tile_97_filtered_output_c11(3);
   bh86_w96_5_c11 <= tile_97_filtered_output_c11(4);
   tile_98_X_c11 <= X(46 downto 44);
   tile_98_Y_c0 <= Y(52 downto 51);
   tile_98_mult: IntMultiplierLUT_3x2_Freq300_uid473
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_98_X_c11,
                 Y => tile_98_Y_c0,
                 R => tile_98_output_c11);

   tile_98_filtered_output_c11 <= unsigned(tile_98_output_c11(4 downto 0));
   bh86_w95_5_c11 <= tile_98_filtered_output_c11(0);
   bh86_w96_6_c11 <= tile_98_filtered_output_c11(1);
   bh86_w97_5_c11 <= tile_98_filtered_output_c11(2);
   bh86_w98_3_c11 <= tile_98_filtered_output_c11(3);
   bh86_w99_4_c11 <= tile_98_filtered_output_c11(4);
   tile_99_X_c11 <= X(49 downto 47);
   tile_99_Y_c0 <= Y(52 downto 51);
   tile_99_mult: IntMultiplierLUT_3x2_Freq300_uid478
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_99_X_c11,
                 Y => tile_99_Y_c0,
                 R => tile_99_output_c11);

   tile_99_filtered_output_c11 <= unsigned(tile_99_output_c11(4 downto 0));
   bh86_w98_4_c11 <= tile_99_filtered_output_c11(0);
   bh86_w99_5_c11 <= tile_99_filtered_output_c11(1);
   bh86_w100_4_c11 <= tile_99_filtered_output_c11(2);
   bh86_w101_5_c11 <= tile_99_filtered_output_c11(3);
   bh86_w102_5_c11 <= tile_99_filtered_output_c11(4);
   tile_100_X_c11 <= X(16 downto 16);
   tile_100_Y_c0 <= Y(48 downto 48);
   tile_100_mult: IntMultiplierLUT_1x1_Freq300_uid483
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_100_X_c11,
                 Y => tile_100_Y_c0,
                 R => tile_100_output_c11);

   tile_100_filtered_output_c11 <= unsigned(tile_100_output_c11(0 downto 0));
   bh86_w64_4_c11 <= tile_100_filtered_output_c11(0);
   tile_101_X_c11 <= X(20 downto 17);
   tile_101_Y_c0 <= Y(48 downto 48);
   tile_101_mult: IntMultiplierLUT_4x1_Freq300_uid485
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_101_X_c11,
                 Y => tile_101_Y_c0,
                 R => tile_101_output_c11);

   tile_101_filtered_output_c11 <= unsigned(tile_101_output_c11(3 downto 0));
   bh86_w65_4_c11 <= tile_101_filtered_output_c11(0);
   bh86_w66_4_c11 <= tile_101_filtered_output_c11(1);
   bh86_w67_4_c11 <= tile_101_filtered_output_c11(2);
   bh86_w68_4_c11 <= tile_101_filtered_output_c11(3);
   tile_102_X_c11 <= X(24 downto 21);
   tile_102_Y_c0 <= Y(48 downto 48);
   tile_102_mult: IntMultiplierLUT_4x1_Freq300_uid487
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_102_X_c11,
                 Y => tile_102_Y_c0,
                 R => tile_102_output_c11);

   tile_102_filtered_output_c11 <= unsigned(tile_102_output_c11(3 downto 0));
   bh86_w69_4_c11 <= tile_102_filtered_output_c11(0);
   bh86_w70_4_c11 <= tile_102_filtered_output_c11(1);
   bh86_w71_4_c11 <= tile_102_filtered_output_c11(2);
   bh86_w72_4_c11 <= tile_102_filtered_output_c11(3);
   tile_103_X_c11 <= X(28 downto 25);
   tile_103_Y_c0 <= Y(48 downto 48);
   tile_103_mult: IntMultiplierLUT_4x1_Freq300_uid489
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_103_X_c11,
                 Y => tile_103_Y_c0,
                 R => tile_103_output_c11);

   tile_103_filtered_output_c11 <= unsigned(tile_103_output_c11(3 downto 0));
   bh86_w73_4_c11 <= tile_103_filtered_output_c11(0);
   bh86_w74_4_c11 <= tile_103_filtered_output_c11(1);
   bh86_w75_4_c11 <= tile_103_filtered_output_c11(2);
   bh86_w76_4_c11 <= tile_103_filtered_output_c11(3);
   tile_104_X_c11 <= X(32 downto 29);
   tile_104_Y_c0 <= Y(48 downto 48);
   tile_104_mult: IntMultiplierLUT_4x1_Freq300_uid491
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_104_X_c11,
                 Y => tile_104_Y_c0,
                 R => tile_104_output_c11);

   tile_104_filtered_output_c11 <= unsigned(tile_104_output_c11(3 downto 0));
   bh86_w77_4_c11 <= tile_104_filtered_output_c11(0);
   bh86_w78_4_c11 <= tile_104_filtered_output_c11(1);
   bh86_w79_4_c11 <= tile_104_filtered_output_c11(2);
   bh86_w80_4_c11 <= tile_104_filtered_output_c11(3);
   tile_105_X_c11 <= X(17 downto 16);
   tile_105_Y_c0 <= Y(50 downto 49);
   tile_105_mult: IntMultiplierLUT_2x2_Freq300_uid493
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_105_X_c11,
                 Y => tile_105_Y_c0,
                 R => tile_105_output_c11);

   tile_105_filtered_output_c11 <= unsigned(tile_105_output_c11(3 downto 0));
   bh86_w65_5_c11 <= tile_105_filtered_output_c11(0);
   bh86_w66_5_c11 <= tile_105_filtered_output_c11(1);
   bh86_w67_5_c11 <= tile_105_filtered_output_c11(2);
   bh86_w68_5_c11 <= tile_105_filtered_output_c11(3);
   tile_106_X_c11 <= X(20 downto 18);
   tile_106_Y_c0 <= Y(50 downto 49);
   tile_106_mult: IntMultiplierLUT_3x2_Freq300_uid498
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_106_X_c11,
                 Y => tile_106_Y_c0,
                 R => tile_106_output_c11);

   tile_106_filtered_output_c11 <= unsigned(tile_106_output_c11(4 downto 0));
   bh86_w67_6_c11 <= tile_106_filtered_output_c11(0);
   bh86_w68_6_c11 <= tile_106_filtered_output_c11(1);
   bh86_w69_5_c11 <= tile_106_filtered_output_c11(2);
   bh86_w70_5_c11 <= tile_106_filtered_output_c11(3);
   bh86_w71_5_c11 <= tile_106_filtered_output_c11(4);
   tile_107_X_c11 <= X(23 downto 21);
   tile_107_Y_c0 <= Y(50 downto 49);
   tile_107_mult: IntMultiplierLUT_3x2_Freq300_uid503
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_107_X_c11,
                 Y => tile_107_Y_c0,
                 R => tile_107_output_c11);

   tile_107_filtered_output_c11 <= unsigned(tile_107_output_c11(4 downto 0));
   bh86_w70_6_c11 <= tile_107_filtered_output_c11(0);
   bh86_w71_6_c11 <= tile_107_filtered_output_c11(1);
   bh86_w72_5_c11 <= tile_107_filtered_output_c11(2);
   bh86_w73_5_c11 <= tile_107_filtered_output_c11(3);
   bh86_w74_5_c11 <= tile_107_filtered_output_c11(4);
   tile_108_X_c11 <= X(26 downto 24);
   tile_108_Y_c0 <= Y(50 downto 49);
   tile_108_mult: IntMultiplierLUT_3x2_Freq300_uid508
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_108_X_c11,
                 Y => tile_108_Y_c0,
                 R => tile_108_output_c11);

   tile_108_filtered_output_c11 <= unsigned(tile_108_output_c11(4 downto 0));
   bh86_w73_6_c11 <= tile_108_filtered_output_c11(0);
   bh86_w74_6_c11 <= tile_108_filtered_output_c11(1);
   bh86_w75_5_c11 <= tile_108_filtered_output_c11(2);
   bh86_w76_5_c11 <= tile_108_filtered_output_c11(3);
   bh86_w77_5_c11 <= tile_108_filtered_output_c11(4);
   tile_109_X_c11 <= X(29 downto 27);
   tile_109_Y_c0 <= Y(50 downto 49);
   tile_109_mult: IntMultiplierLUT_3x2_Freq300_uid513
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_109_X_c11,
                 Y => tile_109_Y_c0,
                 R => tile_109_output_c11);

   tile_109_filtered_output_c11 <= unsigned(tile_109_output_c11(4 downto 0));
   bh86_w76_6_c11 <= tile_109_filtered_output_c11(0);
   bh86_w77_6_c11 <= tile_109_filtered_output_c11(1);
   bh86_w78_5_c11 <= tile_109_filtered_output_c11(2);
   bh86_w79_5_c11 <= tile_109_filtered_output_c11(3);
   bh86_w80_5_c11 <= tile_109_filtered_output_c11(4);
   tile_110_X_c11 <= X(32 downto 30);
   tile_110_Y_c0 <= Y(50 downto 49);
   tile_110_mult: IntMultiplierLUT_3x2_Freq300_uid518
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_110_X_c11,
                 Y => tile_110_Y_c0,
                 R => tile_110_output_c11);

   tile_110_filtered_output_c11 <= unsigned(tile_110_output_c11(4 downto 0));
   bh86_w79_6_c11 <= tile_110_filtered_output_c11(0);
   bh86_w80_6_c11 <= tile_110_filtered_output_c11(1);
   bh86_w81_4_c11 <= tile_110_filtered_output_c11(2);
   bh86_w82_5_c11 <= tile_110_filtered_output_c11(3);
   bh86_w83_5_c11 <= tile_110_filtered_output_c11(4);
   tile_111_X_c11 <= X(17 downto 16);
   tile_111_Y_c0 <= Y(52 downto 51);
   tile_111_mult: IntMultiplierLUT_2x2_Freq300_uid523
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_111_X_c11,
                 Y => tile_111_Y_c0,
                 R => tile_111_output_c11);

   tile_111_filtered_output_c11 <= unsigned(tile_111_output_c11(3 downto 0));
   bh86_w67_7_c11 <= tile_111_filtered_output_c11(0);
   bh86_w68_7_c11 <= tile_111_filtered_output_c11(1);
   bh86_w69_6_c11 <= tile_111_filtered_output_c11(2);
   bh86_w70_7_c11 <= tile_111_filtered_output_c11(3);
   tile_112_X_c11 <= X(20 downto 18);
   tile_112_Y_c0 <= Y(52 downto 51);
   tile_112_mult: IntMultiplierLUT_3x2_Freq300_uid528
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_112_X_c11,
                 Y => tile_112_Y_c0,
                 R => tile_112_output_c11);

   tile_112_filtered_output_c11 <= unsigned(tile_112_output_c11(4 downto 0));
   bh86_w69_7_c11 <= tile_112_filtered_output_c11(0);
   bh86_w70_8_c11 <= tile_112_filtered_output_c11(1);
   bh86_w71_7_c11 <= tile_112_filtered_output_c11(2);
   bh86_w72_6_c11 <= tile_112_filtered_output_c11(3);
   bh86_w73_7_c11 <= tile_112_filtered_output_c11(4);
   tile_113_X_c11 <= X(23 downto 21);
   tile_113_Y_c0 <= Y(52 downto 51);
   tile_113_mult: IntMultiplierLUT_3x2_Freq300_uid533
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_113_X_c11,
                 Y => tile_113_Y_c0,
                 R => tile_113_output_c11);

   tile_113_filtered_output_c11 <= unsigned(tile_113_output_c11(4 downto 0));
   bh86_w72_7_c11 <= tile_113_filtered_output_c11(0);
   bh86_w73_8_c11 <= tile_113_filtered_output_c11(1);
   bh86_w74_7_c11 <= tile_113_filtered_output_c11(2);
   bh86_w75_6_c11 <= tile_113_filtered_output_c11(3);
   bh86_w76_7_c11 <= tile_113_filtered_output_c11(4);
   tile_114_X_c11 <= X(26 downto 24);
   tile_114_Y_c0 <= Y(52 downto 51);
   tile_114_mult: IntMultiplierLUT_3x2_Freq300_uid538
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_114_X_c11,
                 Y => tile_114_Y_c0,
                 R => tile_114_output_c11);

   tile_114_filtered_output_c11 <= unsigned(tile_114_output_c11(4 downto 0));
   bh86_w75_7_c11 <= tile_114_filtered_output_c11(0);
   bh86_w76_8_c11 <= tile_114_filtered_output_c11(1);
   bh86_w77_7_c11 <= tile_114_filtered_output_c11(2);
   bh86_w78_6_c11 <= tile_114_filtered_output_c11(3);
   bh86_w79_7_c11 <= tile_114_filtered_output_c11(4);
   tile_115_X_c11 <= X(29 downto 27);
   tile_115_Y_c0 <= Y(52 downto 51);
   tile_115_mult: IntMultiplierLUT_3x2_Freq300_uid543
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_115_X_c11,
                 Y => tile_115_Y_c0,
                 R => tile_115_output_c11);

   tile_115_filtered_output_c11 <= unsigned(tile_115_output_c11(4 downto 0));
   bh86_w78_7_c11 <= tile_115_filtered_output_c11(0);
   bh86_w79_8_c11 <= tile_115_filtered_output_c11(1);
   bh86_w80_7_c11 <= tile_115_filtered_output_c11(2);
   bh86_w81_5_c11 <= tile_115_filtered_output_c11(3);
   bh86_w82_6_c11 <= tile_115_filtered_output_c11(4);
   tile_116_X_c11 <= X(32 downto 30);
   tile_116_Y_c0 <= Y(52 downto 51);
   tile_116_mult: IntMultiplierLUT_3x2_Freq300_uid548
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_116_X_c11,
                 Y => tile_116_Y_c0,
                 R => tile_116_output_c11);

   tile_116_filtered_output_c11 <= unsigned(tile_116_output_c11(4 downto 0));
   bh86_w81_6_c11 <= tile_116_filtered_output_c11(0);
   bh86_w82_7_c11 <= tile_116_filtered_output_c11(1);
   bh86_w83_6_c11 <= tile_116_filtered_output_c11(2);
   bh86_w84_7_c11 <= tile_116_filtered_output_c11(3);
   bh86_w85_7_c11 <= tile_116_filtered_output_c11(4);
   tile_117_X_c11 <= X(3 downto 0);
   tile_117_Y_c0 <= Y(48 downto 48);
   tile_117_mult: IntMultiplierLUT_4x1_Freq300_uid553
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_117_X_c11,
                 Y => tile_117_Y_c0,
                 R => tile_117_output_c11);

   tile_117_filtered_output_c11 <= unsigned(tile_117_output_c11(3 downto 0));
   bh86_w48_21_c11 <= tile_117_filtered_output_c11(0);
   bh86_w49_20_c11 <= tile_117_filtered_output_c11(1);
   bh86_w50_20_c11 <= tile_117_filtered_output_c11(2);
   bh86_w51_18_c11 <= tile_117_filtered_output_c11(3);
   tile_118_X_c11 <= X(7 downto 4);
   tile_118_Y_c0 <= Y(48 downto 48);
   tile_118_mult: IntMultiplierLUT_4x1_Freq300_uid555
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_118_X_c11,
                 Y => tile_118_Y_c0,
                 R => tile_118_output_c11);

   tile_118_filtered_output_c11 <= unsigned(tile_118_output_c11(3 downto 0));
   bh86_w52_16_c11 <= tile_118_filtered_output_c11(0);
   bh86_w53_15_c11 <= tile_118_filtered_output_c11(1);
   bh86_w54_13_c11 <= tile_118_filtered_output_c11(2);
   bh86_w55_11_c11 <= tile_118_filtered_output_c11(3);
   tile_119_X_c11 <= X(11 downto 8);
   tile_119_Y_c0 <= Y(48 downto 48);
   tile_119_mult: IntMultiplierLUT_4x1_Freq300_uid557
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_119_X_c11,
                 Y => tile_119_Y_c0,
                 R => tile_119_output_c11);

   tile_119_filtered_output_c11 <= unsigned(tile_119_output_c11(3 downto 0));
   bh86_w56_10_c11 <= tile_119_filtered_output_c11(0);
   bh86_w57_10_c11 <= tile_119_filtered_output_c11(1);
   bh86_w58_8_c11 <= tile_119_filtered_output_c11(2);
   bh86_w59_8_c11 <= tile_119_filtered_output_c11(3);
   tile_120_X_c11 <= X(15 downto 12);
   tile_120_Y_c0 <= Y(48 downto 48);
   tile_120_mult: IntMultiplierLUT_4x1_Freq300_uid559
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_120_X_c11,
                 Y => tile_120_Y_c0,
                 R => tile_120_output_c11);

   tile_120_filtered_output_c11 <= unsigned(tile_120_output_c11(3 downto 0));
   bh86_w60_7_c11 <= tile_120_filtered_output_c11(0);
   bh86_w61_6_c11 <= tile_120_filtered_output_c11(1);
   bh86_w62_5_c11 <= tile_120_filtered_output_c11(2);
   bh86_w63_5_c11 <= tile_120_filtered_output_c11(3);
   tile_121_X_c11 <= X(0 downto 0);
   tile_121_Y_c0 <= Y(50 downto 49);
   tile_121_mult: IntMultiplierLUT_1x2_Freq300_uid561
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_121_X_c11,
                 Y => tile_121_Y_c0,
                 R => tile_121_output_c11);

   tile_121_filtered_output_c11 <= unsigned(tile_121_output_c11(1 downto 0));
   bh86_w49_21_c11 <= tile_121_filtered_output_c11(0);
   bh86_w50_21_c11 <= tile_121_filtered_output_c11(1);
   tile_122_X_c11 <= X(3 downto 1);
   tile_122_Y_c0 <= Y(50 downto 49);
   tile_122_mult: IntMultiplierLUT_3x2_Freq300_uid563
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_122_X_c11,
                 Y => tile_122_Y_c0,
                 R => tile_122_output_c11);

   tile_122_filtered_output_c11 <= unsigned(tile_122_output_c11(4 downto 0));
   bh86_w50_22_c11 <= tile_122_filtered_output_c11(0);
   bh86_w51_19_c11 <= tile_122_filtered_output_c11(1);
   bh86_w52_17_c11 <= tile_122_filtered_output_c11(2);
   bh86_w53_16_c11 <= tile_122_filtered_output_c11(3);
   bh86_w54_14_c11 <= tile_122_filtered_output_c11(4);
   tile_123_X_c11 <= X(6 downto 4);
   tile_123_Y_c0 <= Y(50 downto 49);
   tile_123_mult: IntMultiplierLUT_3x2_Freq300_uid568
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_123_X_c11,
                 Y => tile_123_Y_c0,
                 R => tile_123_output_c11);

   tile_123_filtered_output_c11 <= unsigned(tile_123_output_c11(4 downto 0));
   bh86_w53_17_c11 <= tile_123_filtered_output_c11(0);
   bh86_w54_15_c11 <= tile_123_filtered_output_c11(1);
   bh86_w55_12_c11 <= tile_123_filtered_output_c11(2);
   bh86_w56_11_c11 <= tile_123_filtered_output_c11(3);
   bh86_w57_11_c11 <= tile_123_filtered_output_c11(4);
   tile_124_X_c11 <= X(9 downto 7);
   tile_124_Y_c0 <= Y(50 downto 49);
   tile_124_mult: IntMultiplierLUT_3x2_Freq300_uid573
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_124_X_c11,
                 Y => tile_124_Y_c0,
                 R => tile_124_output_c11);

   tile_124_filtered_output_c11 <= unsigned(tile_124_output_c11(4 downto 0));
   bh86_w56_12_c11 <= tile_124_filtered_output_c11(0);
   bh86_w57_12_c11 <= tile_124_filtered_output_c11(1);
   bh86_w58_9_c11 <= tile_124_filtered_output_c11(2);
   bh86_w59_9_c11 <= tile_124_filtered_output_c11(3);
   bh86_w60_8_c11 <= tile_124_filtered_output_c11(4);
   tile_125_X_c11 <= X(12 downto 10);
   tile_125_Y_c0 <= Y(50 downto 49);
   tile_125_mult: IntMultiplierLUT_3x2_Freq300_uid578
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_125_X_c11,
                 Y => tile_125_Y_c0,
                 R => tile_125_output_c11);

   tile_125_filtered_output_c11 <= unsigned(tile_125_output_c11(4 downto 0));
   bh86_w59_10_c11 <= tile_125_filtered_output_c11(0);
   bh86_w60_9_c11 <= tile_125_filtered_output_c11(1);
   bh86_w61_7_c11 <= tile_125_filtered_output_c11(2);
   bh86_w62_6_c11 <= tile_125_filtered_output_c11(3);
   bh86_w63_6_c11 <= tile_125_filtered_output_c11(4);
   tile_126_X_c11 <= X(15 downto 13);
   tile_126_Y_c0 <= Y(50 downto 49);
   tile_126_mult: IntMultiplierLUT_3x2_Freq300_uid583
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_126_X_c11,
                 Y => tile_126_Y_c0,
                 R => tile_126_output_c11);

   tile_126_filtered_output_c11 <= unsigned(tile_126_output_c11(4 downto 0));
   bh86_w62_7_c11 <= tile_126_filtered_output_c11(0);
   bh86_w63_7_c11 <= tile_126_filtered_output_c11(1);
   bh86_w64_5_c11 <= tile_126_filtered_output_c11(2);
   bh86_w65_6_c11 <= tile_126_filtered_output_c11(3);
   bh86_w66_6_c11 <= tile_126_filtered_output_c11(4);
   tile_127_X_c11 <= X(0 downto 0);
   tile_127_Y_c0 <= Y(52 downto 51);
   tile_127_mult: IntMultiplierLUT_1x2_Freq300_uid588
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_127_X_c11,
                 Y => tile_127_Y_c0,
                 R => tile_127_output_c11);

   tile_127_filtered_output_c11 <= unsigned(tile_127_output_c11(1 downto 0));
   bh86_w51_20_c11 <= tile_127_filtered_output_c11(0);
   bh86_w52_18_c11 <= tile_127_filtered_output_c11(1);
   tile_128_X_c11 <= X(3 downto 1);
   tile_128_Y_c0 <= Y(52 downto 51);
   tile_128_mult: IntMultiplierLUT_3x2_Freq300_uid590
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_128_X_c11,
                 Y => tile_128_Y_c0,
                 R => tile_128_output_c11);

   tile_128_filtered_output_c11 <= unsigned(tile_128_output_c11(4 downto 0));
   bh86_w52_19_c11 <= tile_128_filtered_output_c11(0);
   bh86_w53_18_c11 <= tile_128_filtered_output_c11(1);
   bh86_w54_16_c11 <= tile_128_filtered_output_c11(2);
   bh86_w55_13_c11 <= tile_128_filtered_output_c11(3);
   bh86_w56_13_c11 <= tile_128_filtered_output_c11(4);
   tile_129_X_c11 <= X(6 downto 4);
   tile_129_Y_c0 <= Y(52 downto 51);
   tile_129_mult: IntMultiplierLUT_3x2_Freq300_uid595
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_129_X_c11,
                 Y => tile_129_Y_c0,
                 R => tile_129_output_c11);

   tile_129_filtered_output_c11 <= unsigned(tile_129_output_c11(4 downto 0));
   bh86_w55_14_c11 <= tile_129_filtered_output_c11(0);
   bh86_w56_14_c11 <= tile_129_filtered_output_c11(1);
   bh86_w57_13_c11 <= tile_129_filtered_output_c11(2);
   bh86_w58_10_c11 <= tile_129_filtered_output_c11(3);
   bh86_w59_11_c11 <= tile_129_filtered_output_c11(4);
   tile_130_X_c11 <= X(9 downto 7);
   tile_130_Y_c0 <= Y(52 downto 51);
   tile_130_mult: IntMultiplierLUT_3x2_Freq300_uid600
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_130_X_c11,
                 Y => tile_130_Y_c0,
                 R => tile_130_output_c11);

   tile_130_filtered_output_c11 <= unsigned(tile_130_output_c11(4 downto 0));
   bh86_w58_11_c11 <= tile_130_filtered_output_c11(0);
   bh86_w59_12_c11 <= tile_130_filtered_output_c11(1);
   bh86_w60_10_c11 <= tile_130_filtered_output_c11(2);
   bh86_w61_8_c11 <= tile_130_filtered_output_c11(3);
   bh86_w62_8_c11 <= tile_130_filtered_output_c11(4);
   tile_131_X_c11 <= X(12 downto 10);
   tile_131_Y_c0 <= Y(52 downto 51);
   tile_131_mult: IntMultiplierLUT_3x2_Freq300_uid605
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_131_X_c11,
                 Y => tile_131_Y_c0,
                 R => tile_131_output_c11);

   tile_131_filtered_output_c11 <= unsigned(tile_131_output_c11(4 downto 0));
   bh86_w61_9_c11 <= tile_131_filtered_output_c11(0);
   bh86_w62_9_c11 <= tile_131_filtered_output_c11(1);
   bh86_w63_8_c11 <= tile_131_filtered_output_c11(2);
   bh86_w64_6_c11 <= tile_131_filtered_output_c11(3);
   bh86_w65_7_c11 <= tile_131_filtered_output_c11(4);
   tile_132_X_c11 <= X(15 downto 13);
   tile_132_Y_c0 <= Y(52 downto 51);
   tile_132_mult: IntMultiplierLUT_3x2_Freq300_uid610
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => tile_132_X_c11,
                 Y => tile_132_Y_c0,
                 R => tile_132_output_c11);

   tile_132_filtered_output_c11 <= unsigned(tile_132_output_c11(4 downto 0));
   bh86_w64_7_c11 <= tile_132_filtered_output_c11(0);
   bh86_w65_8_c11 <= tile_132_filtered_output_c11(1);
   bh86_w66_7_c11 <= tile_132_filtered_output_c11(2);
   bh86_w67_8_c11 <= tile_132_filtered_output_c11(3);
   bh86_w68_8_c11 <= tile_132_filtered_output_c11(4);

   -- Adding the constant bits 
   bh86_w44_30_c0 <= '1';
   bh86_w45_20_c0 <= '1';
   bh86_w46_20_c0 <= '1';
   bh86_w47_24_c0 <= '1';
   bh86_w48_22_c0 <= '1';
   bh86_w49_22_c0 <= '1';


   Compressor_6_3_Freq300_uid616_bh86_uid617_In0_c11 <= "" & bh86_w44_30_c11 & bh86_w44_14_c11 & bh86_w44_29_c11 & bh86_w44_28_c11 & bh86_w44_27_c11 & bh86_w44_26_c11;
   bh86_w44_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_c12(0);
   bh86_w45_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_c12(1);
   bh86_w46_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid617: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid617_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_copy618_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid617_Out0_copy618_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid619_In0_c11 <= "" & bh86_w44_1_c11 & bh86_w44_2_c11 & bh86_w44_3_c11 & bh86_w44_4_c11 & bh86_w44_5_c11 & bh86_w44_6_c11;
   bh86_w44_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_c12(0);
   bh86_w45_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_c12(1);
   bh86_w46_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid619: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid619_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_copy620_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid619_Out0_copy620_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid621_In0_c11 <= "" & bh86_w44_25_c11 & bh86_w44_24_c11 & bh86_w44_23_c11 & bh86_w44_22_c11 & bh86_w44_21_c11 & bh86_w44_20_c11;
   bh86_w44_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_c12(0);
   bh86_w45_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_c12(1);
   bh86_w46_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid621: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid621_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_copy622_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid621_Out0_copy622_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid623_In0_c11 <= "" & bh86_w44_17_c11 & bh86_w44_7_c11 & bh86_w44_8_c11 & bh86_w44_9_c11 & bh86_w44_10_c11 & bh86_w44_11_c11;
   bh86_w44_34_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_c12(0);
   bh86_w45_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_c12(1);
   bh86_w46_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid623: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid623_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_copy624_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid623_Out0_copy624_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid627_In0_c11 <= "" & bh86_w44_15_c11 & bh86_w44_19_c11 & bh86_w44_18_c11 & bh86_w44_16_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c0 <= "" & bh86_w45_20_c0;
   bh86_w44_35_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_c12(0);
   bh86_w45_25_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_c12(1);
   bh86_w46_25_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid627: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid627_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid627_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_copy628_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid627_Out0_copy628_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid629_In0_c11 <= "" & bh86_w45_6_c11 & bh86_w45_12_c11 & bh86_w45_1_c11 & bh86_w45_2_c11 & bh86_w45_3_c11 & bh86_w45_4_c11;
   bh86_w45_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_c12(0);
   bh86_w46_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_c12(1);
   bh86_w47_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid629: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid629_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_copy630_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid629_Out0_copy630_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid631_In0_c11 <= "" & bh86_w45_14_c11 & bh86_w45_10_c11 & bh86_w45_9_c11 & bh86_w45_19_c11 & bh86_w45_18_c11 & bh86_w45_17_c11;
   bh86_w45_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_c12(0);
   bh86_w46_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_c12(1);
   bh86_w47_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid631: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid631_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_copy632_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid631_Out0_copy632_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid633_In0_c11 <= "" & bh86_w45_5_c11 & bh86_w45_7_c11 & bh86_w45_11_c11 & bh86_w45_15_c11 & bh86_w45_16_c11 & bh86_w45_13_c11;
   bh86_w45_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_c12(0);
   bh86_w46_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_c12(1);
   bh86_w47_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid633: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid633_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_copy634_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid633_Out0_copy634_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid635_In0_c11 <= "" & bh86_w46_20_c11 & bh86_w46_10_c11 & bh86_w46_13_c11 & bh86_w46_16_c11 & bh86_w46_17_c11 & bh86_w46_18_c11;
   bh86_w46_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_c12(0);
   bh86_w47_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_c12(1);
   bh86_w48_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid635: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid635_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_copy636_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid635_Out0_copy636_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid637_In0_c11 <= "" & bh86_w46_2_c11 & bh86_w46_11_c11 & bh86_w46_5_c11 & bh86_w46_6_c11 & bh86_w46_12_c11 & bh86_w46_1_c11;
   bh86_w46_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_c12(0);
   bh86_w47_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_c12(1);
   bh86_w48_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid637: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid637_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_copy638_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid637_Out0_copy638_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid639_In0_c11 <= "" & bh86_w46_15_c11 & bh86_w46_19_c11 & bh86_w46_9_c11 & bh86_w46_14_c11 & bh86_w46_4_c11 & bh86_w46_3_c11;
   bh86_w46_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_c12(0);
   bh86_w47_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_c12(1);
   bh86_w48_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid639: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid639_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_copy640_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid639_Out0_copy640_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid641_In0_c11 <= "" & bh86_w47_24_c11 & bh86_w47_10_c11 & bh86_w47_14_c11 & bh86_w47_11_c11 & "0" & "0";
   bh86_w47_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_c12(0);
   bh86_w48_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_c12(1);
   bh86_w49_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid641: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid641_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_copy642_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid641_Out0_copy642_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid643_In0_c11 <= "" & bh86_w47_15_c11 & bh86_w47_13_c11 & bh86_w47_12_c11 & bh86_w47_23_c11 & bh86_w47_22_c11 & bh86_w47_21_c11;
   bh86_w47_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_c12(0);
   bh86_w48_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_c12(1);
   bh86_w49_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid643: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid643_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_copy644_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid643_Out0_copy644_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid645_In0_c11 <= "" & bh86_w47_8_c11 & bh86_w47_1_c11 & bh86_w47_2_c11 & bh86_w47_3_c11 & bh86_w47_4_c11 & bh86_w47_5_c11;
   bh86_w47_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_c12(0);
   bh86_w48_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_c12(1);
   bh86_w49_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid645: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid645_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_copy646_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid645_Out0_copy646_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid647_In0_c11 <= "" & bh86_w47_17_c11 & bh86_w47_20_c11 & bh86_w47_19_c11 & bh86_w47_18_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c0 <= "" & bh86_w48_22_c0;
   bh86_w47_34_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_c12(0);
   bh86_w48_29_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_c12(1);
   bh86_w49_26_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid647: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid647_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid647_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_copy648_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid647_Out0_copy648_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid651_In0_c11 <= "" & bh86_w47_6_c11 & bh86_w47_7_c11 & bh86_w47_16_c11;
   Compressor_23_3_Freq300_uid650_bh86_uid651_In1_c11 <= "" & bh86_w48_5_c11 & bh86_w48_12_c11;
   bh86_w47_35_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_c12(0);
   bh86_w48_30_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_c12(1);
   bh86_w49_27_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid651: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid651_In0_c11,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid651_In1_c11,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_copy652_c11);
   Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid651_Out0_copy652_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid653_In0_c11 <= "" & bh86_w48_11_c11 & bh86_w48_15_c11 & bh86_w48_17_c11 & bh86_w48_18_c11 & bh86_w48_19_c11 & bh86_w48_20_c11;
   bh86_w48_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_c12(0);
   bh86_w49_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_c12(1);
   bh86_w50_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid653: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid653_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_copy654_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid653_Out0_copy654_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid655_In0_c11 <= "" & bh86_w48_13_c11 & bh86_w48_9_c11 & bh86_w48_6_c11 & bh86_w48_4_c11 & bh86_w48_3_c11 & bh86_w48_2_c11;
   bh86_w48_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_c12(0);
   bh86_w49_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_c12(1);
   bh86_w50_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid655: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid655_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_copy656_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid655_Out0_copy656_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid657_In0_c11 <= "" & bh86_w48_16_c11 & bh86_w48_21_c11 & bh86_w48_10_c11 & bh86_w48_14_c11 & bh86_w48_1_c11 & bh86_w48_7_c11;
   bh86_w48_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_c12(0);
   bh86_w49_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_c12(1);
   bh86_w50_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid657: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid657_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_copy658_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid657_Out0_copy658_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid659_In0_c11 <= "" & bh86_w49_22_c11 & bh86_w49_9_c11 & bh86_w49_12_c11 & bh86_w49_5_c11 & bh86_w49_4_c11 & bh86_w49_3_c11;
   bh86_w49_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_c12(0);
   bh86_w50_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_c12(1);
   bh86_w51_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid659: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid659_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_copy660_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid659_Out0_copy660_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid661_In0_c11 <= "" & bh86_w49_16_c11 & bh86_w49_15_c11 & bh86_w49_21_c11 & bh86_w49_20_c11 & bh86_w49_19_c11 & bh86_w49_18_c11;
   bh86_w49_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_c12(0);
   bh86_w50_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_c12(1);
   bh86_w51_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid661: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid661_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_copy662_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid661_Out0_copy662_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid663_In0_c11 <= "" & bh86_w49_2_c11 & bh86_w49_6_c11 & bh86_w49_1_c11 & bh86_w49_10_c11 & bh86_w49_8_c11 & bh86_w49_11_c11;
   bh86_w49_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_c12(0);
   bh86_w50_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_c12(1);
   bh86_w51_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid663: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid663_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_copy664_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid663_Out0_copy664_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid665_In0_c11 <= "" & bh86_w49_14_c11 & bh86_w49_17_c11 & bh86_w49_13_c11;
   Compressor_23_3_Freq300_uid650_bh86_uid665_In1_c11 <= "" & bh86_w50_22_c11 & bh86_w50_14_c11;
   bh86_w49_34_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_c12(0);
   bh86_w50_29_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_c12(1);
   bh86_w51_24_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid665: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid665_In0_c11,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid665_In1_c11,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_copy666_c11);
   Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid665_Out0_copy666_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid667_In0_c11 <= "" & bh86_w50_12_c11 & bh86_w50_11_c11 & bh86_w50_3_c11 & bh86_w50_4_c11 & bh86_w50_5_c11 & bh86_w50_6_c11;
   bh86_w50_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_c12(0);
   bh86_w51_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_c12(1);
   bh86_w52_20_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid667: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid667_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_copy668_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid667_Out0_copy668_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid669_In0_c11 <= "" & bh86_w50_15_c11 & bh86_w50_16_c11 & bh86_w50_17_c11 & bh86_w50_18_c11 & bh86_w50_19_c11 & bh86_w50_20_c11;
   bh86_w50_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_c12(0);
   bh86_w51_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_c12(1);
   bh86_w52_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid669: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid669_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_copy670_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid669_Out0_copy670_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid671_In0_c11 <= "" & bh86_w50_10_c11 & bh86_w50_7_c11 & bh86_w50_9_c11 & bh86_w50_13_c11 & bh86_w50_21_c11 & bh86_w50_2_c11;
   bh86_w50_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_c12(0);
   bh86_w51_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_c12(1);
   bh86_w52_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid671: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid671_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_copy672_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid671_Out0_copy672_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid673_In0_c11 <= "" & bh86_w51_20_c11 & bh86_w51_13_c11 & bh86_w51_10_c11 & bh86_w51_19_c11 & bh86_w51_18_c11 & bh86_w51_17_c11;
   bh86_w51_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_c12(0);
   bh86_w52_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_c12(1);
   bh86_w53_19_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid673: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid673_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_copy674_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid673_Out0_copy674_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid675_In0_c11 <= "" & bh86_w51_11_c11 & bh86_w51_2_c11 & bh86_w51_3_c11 & bh86_w51_4_c11 & bh86_w51_5_c11 & bh86_w51_7_c11;
   bh86_w51_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_c12(0);
   bh86_w52_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_c12(1);
   bh86_w53_20_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid675: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid675_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_copy676_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid675_Out0_copy676_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid677_In0_c11 <= "" & bh86_w51_14_c11 & bh86_w51_16_c11 & bh86_w51_15_c11 & bh86_w51_12_c11 & bh86_w51_8_c11 & bh86_w51_9_c11;
   bh86_w51_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_c12(0);
   bh86_w52_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_c12(1);
   bh86_w53_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid677: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid677_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_copy678_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid677_Out0_copy678_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid679_In0_c11 <= "" & bh86_w52_2_c11 & bh86_w52_10_c11 & bh86_w52_3_c11 & bh86_w52_4_c11 & bh86_w52_5_c11 & bh86_w52_7_c11;
   bh86_w52_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_c12(0);
   bh86_w53_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_c12(1);
   bh86_w54_17_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid679: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid679_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_copy680_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid679_Out0_copy680_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid681_In0_c11 <= "" & bh86_w52_12_c11 & bh86_w52_19_c11 & bh86_w52_18_c11 & bh86_w52_17_c11 & bh86_w52_16_c11 & bh86_w52_15_c11;
   bh86_w52_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_c12(0);
   bh86_w53_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_c12(1);
   bh86_w54_18_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid681: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid681_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_copy682_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid681_Out0_copy682_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid683_In0_c11 <= "" & bh86_w52_11_c11 & bh86_w52_8_c11 & bh86_w52_9_c11 & bh86_w52_14_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid683_In1_c11 <= "" & bh86_w53_2_c11;
   bh86_w52_28_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_c12(0);
   bh86_w53_24_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_c12(1);
   bh86_w54_19_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid683: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid683_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid683_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_copy684_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid683_Out0_copy684_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid685_In0_c11 <= "" & bh86_w53_9_c11 & bh86_w53_17_c11 & bh86_w53_16_c11 & bh86_w53_15_c11 & bh86_w53_14_c11 & bh86_w53_13_c11;
   bh86_w53_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_c12(0);
   bh86_w54_20_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_c12(1);
   bh86_w55_15_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid685: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid685_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_copy686_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid685_Out0_copy686_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid687_In0_c11 <= "" & bh86_w53_18_c11 & bh86_w53_3_c11 & bh86_w53_4_c11 & bh86_w53_6_c11 & bh86_w53_7_c11 & bh86_w53_8_c11;
   bh86_w53_26_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_c12(0);
   bh86_w54_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_c12(1);
   bh86_w55_16_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid687: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid687_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_copy688_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid687_Out0_copy688_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid689_In0_c11 <= "" & bh86_w53_12_c11 & bh86_w53_11_c11 & bh86_w53_10_c11;
   Compressor_23_3_Freq300_uid650_bh86_uid689_In1_c11 <= "" & bh86_w54_2_c11 & bh86_w54_16_c11;
   bh86_w53_27_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_c12(0);
   bh86_w54_22_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_c12(1);
   bh86_w55_17_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid689: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid689_In0_c11,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid689_In1_c11,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_copy690_c11);
   Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid689_Out0_copy690_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid691_In0_c11 <= "" & bh86_w54_8_c11 & bh86_w54_3_c11 & bh86_w54_5_c11 & bh86_w54_6_c11 & bh86_w54_7_c11 & bh86_w54_9_c11;
   bh86_w54_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_c12(0);
   bh86_w55_18_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_c12(1);
   bh86_w56_15_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid691: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid691_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_copy692_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid691_Out0_copy692_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid693_In0_c11 <= "" & bh86_w54_15_c11 & bh86_w54_14_c11 & bh86_w54_13_c11 & bh86_w54_12_c11 & bh86_w54_11_c11 & bh86_w54_10_c11;
   bh86_w54_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_c12(0);
   bh86_w55_19_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_c12(1);
   bh86_w56_16_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid693: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid693_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_copy694_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid693_Out0_copy694_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid695_In0_c11 <= "" & bh86_w55_2_c11 & bh86_w55_4_c11 & bh86_w55_5_c11 & bh86_w55_6_c11 & bh86_w55_7_c11 & bh86_w55_8_c11;
   bh86_w55_20_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_c12(0);
   bh86_w56_17_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_c12(1);
   bh86_w57_14_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid695: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid695_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_copy696_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid695_Out0_copy696_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid697_In0_c11 <= "" & bh86_w55_14_c11 & bh86_w55_13_c11 & bh86_w55_12_c11 & bh86_w55_11_c11 & bh86_w55_10_c11 & bh86_w55_9_c11;
   bh86_w55_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_c12(0);
   bh86_w56_18_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_c12(1);
   bh86_w57_15_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid697: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid697_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_copy698_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid697_Out0_copy698_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid699_In0_c11 <= "" & bh86_w56_2_c11 & bh86_w56_14_c11 & bh86_w56_13_c11 & bh86_w56_12_c11 & bh86_w56_11_c11 & bh86_w56_10_c11;
   bh86_w56_19_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_c12(0);
   bh86_w57_16_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_c12(1);
   bh86_w58_12_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid699: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid699_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_copy700_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid699_Out0_copy700_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid701_In0_c11 <= "" & bh86_w56_4_c11 & bh86_w56_5_c11 & bh86_w56_6_c11 & bh86_w56_7_c11 & bh86_w56_8_c11 & bh86_w56_9_c11;
   bh86_w56_20_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_c12(0);
   bh86_w57_17_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_c12(1);
   bh86_w58_13_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid701: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid701_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_copy702_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid701_Out0_copy702_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid703_In0_c11 <= "" & bh86_w57_4_c11 & bh86_w57_5_c11 & bh86_w57_6_c11 & bh86_w57_7_c11 & bh86_w57_8_c11 & bh86_w57_9_c11;
   bh86_w57_18_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_c12(0);
   bh86_w58_14_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_c12(1);
   bh86_w59_13_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid703: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid703_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_copy704_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid703_Out0_copy704_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid705_In0_c11 <= "" & bh86_w57_13_c11 & bh86_w57_12_c11 & bh86_w57_11_c11 & bh86_w57_10_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid705_In1_c11 <= "" & bh86_w58_4_c11;
   bh86_w57_19_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_c12(0);
   bh86_w58_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_c12(1);
   bh86_w59_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid705: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid705_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid705_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_copy706_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid705_Out0_copy706_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid707_In0_c11 <= "" & bh86_w58_5_c11 & bh86_w58_6_c11 & bh86_w58_7_c11 & bh86_w58_8_c11 & bh86_w58_9_c11 & bh86_w58_10_c11;
   bh86_w58_16_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_c12(0);
   bh86_w59_15_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_c12(1);
   bh86_w60_11_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid707: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid707_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_copy708_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid707_Out0_copy708_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid709_In0_c11 <= "" & bh86_w59_4_c11 & bh86_w59_5_c11 & bh86_w59_6_c11 & bh86_w59_7_c11 & bh86_w59_8_c11 & bh86_w59_9_c11;
   bh86_w59_16_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_c12(0);
   bh86_w60_12_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_c12(1);
   bh86_w61_10_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid709: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid709_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_copy710_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid709_Out0_copy710_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid713_In0_c11 <= "" & bh86_w59_12_c11 & bh86_w59_11_c11 & bh86_w59_10_c11;
   bh86_w59_17_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_c12(0);
   bh86_w60_13_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid713: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid713_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_copy714_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid713_Out0_copy714_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid715_In0_c11 <= "" & bh86_w60_4_c11 & bh86_w60_5_c11 & bh86_w60_6_c11 & bh86_w60_7_c11 & bh86_w60_8_c11 & bh86_w60_9_c11;
   bh86_w60_14_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_c12(0);
   bh86_w61_11_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_c12(1);
   bh86_w62_10_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid715: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid715_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_copy716_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid715_Out0_copy716_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid717_In0_c11 <= "" & bh86_w61_4_c11 & bh86_w61_5_c11 & bh86_w61_6_c11 & bh86_w61_7_c11 & bh86_w61_8_c11 & bh86_w61_9_c11;
   bh86_w61_12_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_c12(0);
   bh86_w62_11_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_c12(1);
   bh86_w63_9_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid717: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid717_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_copy718_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid717_Out0_copy718_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid719_In0_c11 <= "" & bh86_w62_4_c11 & bh86_w62_5_c11 & bh86_w62_6_c11 & bh86_w62_7_c11 & bh86_w62_8_c11 & bh86_w62_9_c11;
   bh86_w62_12_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_c12(0);
   bh86_w63_10_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_c12(1);
   bh86_w64_8_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid719: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid719_In0_c11,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_copy720_c11);
   Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid719_Out0_copy720_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid721_In0_c11 <= "" & bh86_w63_4_c11 & bh86_w63_5_c11 & bh86_w63_6_c11 & bh86_w63_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid721_In1_c11 <= "" & bh86_w64_4_c11;
   bh86_w63_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_c12(0);
   bh86_w64_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_c12(1);
   bh86_w65_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid721: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid721_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid721_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_copy722_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid721_Out0_copy722_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid723_In0_c11 <= "" & bh86_w64_5_c11 & bh86_w64_6_c11 & bh86_w64_7_c11;
   bh86_w64_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_c12(0);
   bh86_w65_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid723: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid723_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_copy724_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid723_Out0_copy724_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid725_In0_c11 <= "" & bh86_w65_4_c11 & bh86_w65_5_c11 & bh86_w65_6_c11 & bh86_w65_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid725_In1_c11 <= "" & bh86_w66_4_c11;
   bh86_w65_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_c12(0);
   bh86_w66_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_c12(1);
   bh86_w67_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid725: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid725_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid725_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_copy726_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid725_Out0_copy726_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid727_In0_c11 <= "" & bh86_w66_5_c11 & bh86_w66_6_c11 & bh86_w66_7_c11;
   bh86_w66_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_c12(0);
   bh86_w67_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid727: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid727_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_copy728_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid727_Out0_copy728_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid729_In0_c11 <= "" & bh86_w67_4_c11 & bh86_w67_5_c11 & bh86_w67_6_c11 & bh86_w67_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid729_In1_c11 <= "" & bh86_w68_4_c11;
   bh86_w67_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_c12(0);
   bh86_w68_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_c12(1);
   bh86_w69_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid729: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid729_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid729_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_copy730_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid729_Out0_copy730_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid731_In0_c11 <= "" & bh86_w68_5_c11 & bh86_w68_6_c11 & bh86_w68_7_c11 & bh86_w68_8_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid731_In1_c11 <= "" & bh86_w69_4_c11;
   bh86_w68_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_c12(0);
   bh86_w69_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_c12(1);
   bh86_w70_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid731: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid731_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid731_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_copy732_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid731_Out0_copy732_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid733_In0_c11 <= "" & bh86_w69_5_c11 & bh86_w69_6_c11 & bh86_w69_7_c11;
   bh86_w69_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_c12(0);
   bh86_w70_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid733: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid733_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_copy734_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid733_Out0_copy734_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid735_In0_c11 <= "" & bh86_w70_4_c11 & bh86_w70_5_c11 & bh86_w70_6_c11 & bh86_w70_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid735_In1_c11 <= "" & bh86_w71_4_c11;
   bh86_w70_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_c12(0);
   bh86_w71_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_c12(1);
   bh86_w72_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid735: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid735_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid735_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_copy736_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid735_Out0_copy736_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid737_In0_c11 <= "" & bh86_w71_5_c11 & bh86_w71_6_c11 & bh86_w71_7_c11;
   bh86_w71_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_c12(0);
   bh86_w72_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid737: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid737_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_copy738_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid737_Out0_copy738_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid739_In0_c11 <= "" & bh86_w72_4_c11 & bh86_w72_5_c11 & bh86_w72_6_c11 & bh86_w72_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid739_In1_c11 <= "" & bh86_w73_4_c11;
   bh86_w72_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_c12(0);
   bh86_w73_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_c12(1);
   bh86_w74_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid739: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid739_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid739_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_copy740_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid739_Out0_copy740_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid741_In0_c11 <= "" & bh86_w73_5_c11 & bh86_w73_6_c11 & bh86_w73_7_c11 & bh86_w73_8_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid741_In1_c11 <= "" & bh86_w74_4_c11;
   bh86_w73_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_c12(0);
   bh86_w74_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_c12(1);
   bh86_w75_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid741: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid741_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid741_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_copy742_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid741_Out0_copy742_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid743_In0_c11 <= "" & bh86_w74_5_c11 & bh86_w74_6_c11 & bh86_w74_7_c11;
   bh86_w74_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_c12(0);
   bh86_w75_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid743: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid743_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_copy744_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid743_Out0_copy744_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid745_In0_c11 <= "" & bh86_w75_4_c11 & bh86_w75_5_c11 & bh86_w75_6_c11 & bh86_w75_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid745_In1_c11 <= "" & bh86_w76_4_c11;
   bh86_w75_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_c12(0);
   bh86_w76_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_c12(1);
   bh86_w77_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid745: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid745_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid745_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_copy746_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid745_Out0_copy746_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid747_In0_c11 <= "" & bh86_w76_5_c11 & bh86_w76_6_c11 & bh86_w76_7_c11 & bh86_w76_8_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid747_In1_c11 <= "" & bh86_w77_4_c11;
   bh86_w76_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_c12(0);
   bh86_w77_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_c12(1);
   bh86_w78_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid747: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid747_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid747_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_copy748_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid747_Out0_copy748_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid749_In0_c11 <= "" & bh86_w77_5_c11 & bh86_w77_6_c11 & bh86_w77_7_c11;
   bh86_w77_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_c12(0);
   bh86_w78_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid749: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid749_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_copy750_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid749_Out0_copy750_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid751_In0_c11 <= "" & bh86_w78_4_c11 & bh86_w78_5_c11 & bh86_w78_6_c11 & bh86_w78_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid751_In1_c11 <= "" & bh86_w79_4_c11;
   bh86_w78_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_c12(0);
   bh86_w79_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_c12(1);
   bh86_w80_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid751: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid751_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid751_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_copy752_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid751_Out0_copy752_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid753_In0_c11 <= "" & bh86_w79_5_c11 & bh86_w79_6_c11 & bh86_w79_7_c11 & bh86_w79_8_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid753_In1_c11 <= "" & bh86_w80_4_c11;
   bh86_w79_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_c12(0);
   bh86_w80_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_c12(1);
   bh86_w81_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid753: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid753_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid753_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_copy754_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid753_Out0_copy754_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid755_In0_c11 <= "" & bh86_w80_5_c11 & bh86_w80_6_c11 & bh86_w80_7_c11;
   bh86_w80_10_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_c12(0);
   bh86_w81_8_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid755: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid755_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_copy756_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid755_Out0_copy756_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid757_In0_c11 <= "" & bh86_w81_3_c11 & bh86_w81_4_c11 & bh86_w81_5_c11 & bh86_w81_6_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid757_In1_c11 <= "" & bh86_w82_3_c11;
   bh86_w81_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_c12(0);
   bh86_w82_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_c12(1);
   bh86_w83_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid757: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid757_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid757_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_copy758_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid757_Out0_copy758_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid759_In0_c11 <= "" & bh86_w82_4_c11 & bh86_w82_5_c11 & bh86_w82_6_c11 & bh86_w82_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid759_In1_c11 <= "" & bh86_w83_3_c11;
   bh86_w82_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_c12(0);
   bh86_w83_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_c12(1);
   bh86_w84_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid759: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid759_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid759_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_copy760_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid759_Out0_copy760_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid761_In0_c11 <= "" & bh86_w83_4_c11 & bh86_w83_5_c11 & bh86_w83_6_c11;
   bh86_w83_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_c12(0);
   bh86_w84_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid761: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid761_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_copy762_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid761_Out0_copy762_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid763_In0_c11 <= "" & bh86_w84_3_c11 & bh86_w84_4_c11 & bh86_w84_5_c11 & bh86_w84_6_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid763_In1_c11 <= "" & bh86_w85_3_c11;
   bh86_w84_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_c12(0);
   bh86_w85_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_c12(1);
   bh86_w86_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid763: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid763_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid763_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_copy764_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid763_Out0_copy764_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid765_In0_c11 <= "" & bh86_w85_4_c11 & bh86_w85_5_c11 & bh86_w85_6_c11 & bh86_w85_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid765_In1_c11 <= "" & bh86_w86_3_c11;
   bh86_w85_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_c12(0);
   bh86_w86_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_c12(1);
   bh86_w87_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid765: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid765_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid765_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_copy766_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid765_Out0_copy766_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid767_In0_c11 <= "" & bh86_w86_4_c11 & bh86_w86_5_c11 & bh86_w86_6_c11;
   bh86_w86_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_c12(0);
   bh86_w87_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid767: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid767_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_copy768_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid767_Out0_copy768_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid769_In0_c11 <= "" & bh86_w87_3_c11 & bh86_w87_4_c11 & bh86_w87_5_c11 & bh86_w87_6_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid769_In1_c11 <= "" & bh86_w88_3_c11;
   bh86_w87_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_c12(0);
   bh86_w88_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_c12(1);
   bh86_w89_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid769: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid769_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid769_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_copy770_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid769_Out0_copy770_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid771_In0_c11 <= "" & bh86_w88_4_c11 & bh86_w88_5_c11 & bh86_w88_6_c11;
   bh86_w88_8_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_c12(0);
   bh86_w89_8_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid771: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid771_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_copy772_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid771_Out0_copy772_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid773_In0_c11 <= "" & bh86_w89_3_c11 & bh86_w89_4_c11 & bh86_w89_5_c11 & bh86_w89_6_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid773_In1_c11 <= "" & bh86_w90_3_c11;
   bh86_w89_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_c12(0);
   bh86_w90_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_c12(1);
   bh86_w91_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid773: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid773_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid773_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_copy774_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid773_Out0_copy774_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid775_In0_c11 <= "" & bh86_w90_4_c11 & bh86_w90_5_c11 & bh86_w90_6_c11 & bh86_w90_7_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid775_In1_c11 <= "" & bh86_w91_2_c11;
   bh86_w90_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_c12(0);
   bh86_w91_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_c12(1);
   bh86_w92_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid775: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid775_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid775_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_copy776_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid775_Out0_copy776_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid777_In0_c11 <= "" & bh86_w91_3_c11 & bh86_w91_4_c11 & bh86_w91_5_c11;
   bh86_w91_8_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_c12(0);
   bh86_w92_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid777: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid777_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_copy778_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid777_Out0_copy778_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid779_In0_c11 <= "" & bh86_w92_2_c11 & bh86_w92_3_c11 & bh86_w92_4_c11 & bh86_w92_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid779_In1_c11 <= "" & bh86_w93_2_c11;
   bh86_w92_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_c12(0);
   bh86_w93_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_c12(1);
   bh86_w94_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid779: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid779_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid779_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_copy780_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid779_Out0_copy780_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid781_In0_c11 <= "" & bh86_w93_3_c11 & bh86_w93_4_c11 & bh86_w93_5_c11 & bh86_w93_6_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid781_In1_c11 <= "" & bh86_w94_2_c11;
   bh86_w93_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_c12(0);
   bh86_w94_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_c12(1);
   bh86_w95_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid781: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid781_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid781_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_copy782_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid781_Out0_copy782_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid783_In0_c11 <= "" & bh86_w94_3_c11 & bh86_w94_4_c11 & bh86_w94_5_c11;
   bh86_w94_8_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_c12(0);
   bh86_w95_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid783: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid783_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_copy784_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid783_Out0_copy784_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid785_In0_c11 <= "" & bh86_w95_2_c11 & bh86_w95_3_c11 & bh86_w95_4_c11 & bh86_w95_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid785_In1_c11 <= "" & bh86_w96_2_c11;
   bh86_w95_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_c12(0);
   bh86_w96_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_c12(1);
   bh86_w97_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid785: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid785_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid785_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_copy786_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid785_Out0_copy786_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid787_In0_c11 <= "" & bh86_w96_3_c11 & bh86_w96_4_c11 & bh86_w96_5_c11 & bh86_w96_6_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid787_In1_c11 <= "" & bh86_w97_2_c11;
   bh86_w96_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_c12(0);
   bh86_w97_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_c12(1);
   bh86_w98_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid787: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid787_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid787_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_copy788_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid787_Out0_copy788_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid789_In0_c11 <= "" & bh86_w97_3_c11 & bh86_w97_4_c11 & bh86_w97_5_c11;
   bh86_w97_8_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_c12(0);
   bh86_w98_6_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid789: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid789_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_copy790_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid789_Out0_copy790_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid791_In0_c11 <= "" & bh86_w98_1_c11 & bh86_w98_2_c11 & bh86_w98_3_c11 & bh86_w98_4_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid791_In1_c11 <= "" & bh86_w99_1_c11;
   bh86_w98_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_c12(0);
   bh86_w99_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_c12(1);
   bh86_w100_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid791: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid791_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid791_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_copy792_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid791_Out0_copy792_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid793_In0_c11 <= "" & bh86_w99_2_c11 & bh86_w99_3_c11 & bh86_w99_4_c11 & bh86_w99_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid793_In1_c11 <= "" & bh86_w100_1_c11;
   bh86_w99_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_c12(0);
   bh86_w100_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_c12(1);
   bh86_w101_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid793: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid793_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid793_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_copy794_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid793_Out0_copy794_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid795_In0_c11 <= "" & bh86_w100_2_c11 & bh86_w100_3_c11 & bh86_w100_4_c11;
   bh86_w100_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_c12(0);
   bh86_w101_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid795: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid795_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_copy796_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid795_Out0_copy796_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid797_In0_c11 <= "" & bh86_w101_1_c11 & bh86_w101_2_c11 & bh86_w101_3_c11 & bh86_w101_4_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid797_In1_c11 <= "" & bh86_w102_1_c11;
   bh86_w101_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_c12(0);
   bh86_w102_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_c12(1);
   bh86_w103_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid797: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid797_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid797_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_copy798_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid797_Out0_copy798_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid799_In0_c11 <= "" & bh86_w102_2_c11 & bh86_w102_3_c11 & bh86_w102_4_c11 & bh86_w102_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid799_In1_c11 <= "" & bh86_w103_1_c11;
   bh86_w102_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_c12(0);
   bh86_w103_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_c12(1);
   bh86_w104_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid799: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid799_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid799_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_copy800_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid799_Out0_copy800_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid801_In0_c11 <= "" & bh86_w103_2_c11 & bh86_w103_3_c11 & bh86_w103_4_c11;
   bh86_w103_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_c12(0);
   bh86_w104_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid801: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid801_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_copy802_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid801_Out0_copy802_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid803_In0_c11 <= "" & bh86_w104_1_c11 & bh86_w104_2_c11 & bh86_w104_3_c11 & bh86_w104_4_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid803_In1_c11 <= "" & bh86_w105_1_c11;
   bh86_w104_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_c12(0);
   bh86_w105_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_c12(1);
   bh86_w106_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid803: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid803_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid803_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_copy804_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid803_Out0_copy804_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid805_In0_c11 <= "" & bh86_w105_2_c11 & bh86_w105_3_c11 & bh86_w105_4_c11;
   bh86_w105_6_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_c12(0);
   bh86_w106_6_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid805: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid805_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_copy806_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid805_Out0_copy806_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid807_In0_c11 <= "" & bh86_w106_1_c11 & bh86_w106_2_c11 & bh86_w106_3_c11 & bh86_w106_4_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid807_In1_c11 <= "" & bh86_w107_1_c11;
   bh86_w106_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_c12(0);
   bh86_w107_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_c12(1);
   bh86_w108_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid807: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid807_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid807_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_copy808_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid807_Out0_copy808_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid809_In0_c11 <= "" & bh86_w107_2_c11 & bh86_w107_3_c11 & bh86_w107_4_c11 & bh86_w107_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid809_In1_c11 <= "" & bh86_w108_1_c11;
   bh86_w107_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_c12(0);
   bh86_w108_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_c12(1);
   bh86_w109_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid809: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid809_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid809_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_copy810_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid809_Out0_copy810_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid811_In0_c11 <= "" & bh86_w108_2_c11 & bh86_w108_3_c11 & bh86_w108_4_c11;
   bh86_w108_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_c12(0);
   bh86_w109_6_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid811: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid811_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_copy812_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid811_Out0_copy812_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid813_In0_c11 <= "" & bh86_w109_1_c11 & bh86_w109_2_c11 & bh86_w109_3_c11 & bh86_w109_4_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid813_In1_c11 <= "" & bh86_w110_1_c11;
   bh86_w109_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_c12(0);
   bh86_w110_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_c12(1);
   bh86_w111_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid813: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid813_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid813_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_copy814_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid813_Out0_copy814_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid815_In0_c11 <= "" & bh86_w110_2_c11 & bh86_w110_3_c11 & bh86_w110_4_c11 & bh86_w110_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid815_In1_c11 <= "" & bh86_w111_1_c11;
   bh86_w110_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_c12(0);
   bh86_w111_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_c12(1);
   bh86_w112_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid815: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid815_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid815_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_copy816_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid815_Out0_copy816_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid817_In0_c11 <= "" & bh86_w111_2_c11 & bh86_w111_3_c11 & bh86_w111_4_c11;
   bh86_w111_7_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_c12(0);
   bh86_w112_6_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid817: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid817_In0_c11,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_copy818_c11);
   Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid817_Out0_copy818_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid819_In0_c11 <= "" & bh86_w112_1_c11 & bh86_w112_2_c11 & bh86_w112_3_c11 & bh86_w112_4_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid819_In1_c11 <= "" & bh86_w113_1_c11;
   bh86_w112_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_c12(0);
   bh86_w113_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_c12(1);
   bh86_w114_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid819: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid819_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid819_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_copy820_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid819_Out0_copy820_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid821_In0_c11 <= "" & bh86_w113_2_c11 & bh86_w113_3_c11 & bh86_w113_4_c11 & bh86_w113_5_c11;
   Compressor_14_3_Freq300_uid626_bh86_uid821_In1_c11 <= "" & bh86_w114_1_c11;
   bh86_w113_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_c12(0);
   bh86_w114_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_c12(1);
   bh86_w115_3_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid821: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid821_In0_c11,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid821_In1_c11,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_copy822_c11);
   Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid821_Out0_copy822_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid823_In0_c11 <= "" & bh86_w114_2_c11 & bh86_w114_3_c11 & bh86_w114_4_c11;
   Compressor_23_3_Freq300_uid650_bh86_uid823_In1_c11 <= "" & bh86_w115_0_c11 & bh86_w115_1_c11;
   bh86_w114_7_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_c12(0);
   bh86_w115_4_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_c12(1);
   bh86_w116_3_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid823: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid823_In0_c11,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid823_In1_c11,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_copy824_c11);
   Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid823_Out0_copy824_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid825_In0_c11 <= "" & bh86_w116_0_c11 & bh86_w116_1_c11 & bh86_w116_2_c11;
   Compressor_23_3_Freq300_uid650_bh86_uid825_In1_c11 <= "" & bh86_w117_0_c11 & bh86_w117_1_c11;
   bh86_w116_4_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_c12(0);
   bh86_w117_2_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_c12(1);
   bh86_w118_1_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid825: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid825_In0_c11,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid825_In1_c11,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_copy826_c11);
   Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid825_Out0_copy826_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid827_In0_c12 <= "" & bh86_w44_35_c12 & bh86_w44_12_c12 & bh86_w44_34_c12 & bh86_w44_32_c12 & bh86_w44_31_c12 & bh86_w44_33_c12;
   bh86_w44_36_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_c12(0);
   bh86_w45_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_c12(1);
   bh86_w46_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid827: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid827_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_copy828_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid827_Out0_copy828_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid829_In0_c12 <= "" & bh86_w45_25_c12 & bh86_w45_28_c12 & bh86_w45_23_c12 & bh86_w45_21_c12 & bh86_w45_22_c12 & "0";
   bh86_w45_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_c12(0);
   bh86_w46_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_c12(1);
   bh86_w47_36_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid829: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid829_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_copy830_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid829_Out0_copy830_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid831_In0_c12 <= "" & bh86_w45_24_c12 & bh86_w45_26_c12 & bh86_w45_27_c12;
   bh86_w45_31_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_c12(0);
   bh86_w46_34_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid831: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid831_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_copy832_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid831_Out0_copy832_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid833_In0_c12 <= "" & bh86_w46_25_c12 & bh86_w46_7_c12 & bh86_w46_23_c12 & bh86_w46_29_c12 & bh86_w46_27_c12 & bh86_w46_26_c12;
   bh86_w46_35_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_c12(0);
   bh86_w47_37_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_c12(1);
   bh86_w48_34_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid833: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid833_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_copy834_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid833_Out0_copy834_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid835_In0_c12 <= "" & bh86_w46_24_c12 & bh86_w46_30_c12 & bh86_w46_31_c12 & bh86_w46_28_c12 & bh86_w46_21_c12 & bh86_w46_22_c12;
   bh86_w46_36_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_c12(0);
   bh86_w47_38_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_c12(1);
   bh86_w48_35_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid835: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid835_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_copy836_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid835_Out0_copy836_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid837_In0_c12 <= "" & bh86_w47_34_c12 & bh86_w47_35_c12 & bh86_w47_33_c12 & bh86_w47_32_c12 & bh86_w47_30_c12 & bh86_w47_28_c12;
   bh86_w47_39_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_c12(0);
   bh86_w48_36_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_c12(1);
   bh86_w49_35_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid837: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid837_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_copy838_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid837_Out0_copy838_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid839_In0_c12 <= "" & bh86_w47_31_c12 & bh86_w47_29_c12 & bh86_w47_27_c12 & bh86_w47_25_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid839_In1_c12 <= "" & bh86_w48_29_c12;
   bh86_w47_40_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_c12(0);
   bh86_w48_37_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_c12(1);
   bh86_w49_36_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid839: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid839_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid839_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_copy840_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid839_Out0_copy840_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid841_In0_c12 <= "" & bh86_w48_30_c12 & bh86_w48_25_c12 & bh86_w48_32_c12 & bh86_w48_28_c12 & bh86_w48_26_c12 & bh86_w48_24_c12;
   bh86_w48_38_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_c12(0);
   bh86_w49_37_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_c12(1);
   bh86_w50_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid841: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid841_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_copy842_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid841_Out0_copy842_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid843_In0_c12 <= "" & bh86_w48_33_c12 & bh86_w48_31_c12 & bh86_w48_27_c12;
   bh86_w48_39_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_c12(0);
   bh86_w49_38_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid843: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid843_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_copy844_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid843_Out0_copy844_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid845_In0_c12 <= "" & bh86_w49_26_c12 & bh86_w49_34_c12 & bh86_w49_27_c12 & bh86_w49_23_c12 & bh86_w49_33_c12 & bh86_w49_32_c12;
   bh86_w49_39_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_c12(0);
   bh86_w50_34_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_c12(1);
   bh86_w51_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid845: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid845_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_copy846_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid845_Out0_copy846_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid847_In0_c12 <= "" & bh86_w49_29_c12 & bh86_w49_30_c12 & bh86_w49_31_c12 & bh86_w49_24_c12 & bh86_w49_25_c12 & bh86_w49_28_c12;
   bh86_w49_40_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_c12(0);
   bh86_w50_35_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_c12(1);
   bh86_w51_32_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid847: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid847_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_copy848_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid847_Out0_copy848_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid849_In0_c12 <= "" & bh86_w50_29_c12 & bh86_w50_31_c12 & bh86_w50_27_c12 & bh86_w50_26_c12 & bh86_w50_25_c12 & bh86_w50_24_c12;
   bh86_w50_36_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_c12(0);
   bh86_w51_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_c12(1);
   bh86_w52_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid849: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid849_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_copy850_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid849_Out0_copy850_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid851_In0_c12 <= "" & bh86_w50_23_c12 & bh86_w50_28_c12 & bh86_w50_30_c12 & bh86_w50_32_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid851_In1_c12 <= "" & bh86_w51_24_c12;
   bh86_w50_37_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_c12(0);
   bh86_w51_34_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_c12(1);
   bh86_w52_30_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid851: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid851_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid851_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_copy852_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid851_Out0_copy852_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid853_In0_c12 <= "" & bh86_w51_29_c12 & bh86_w51_30_c12 & bh86_w51_25_c12 & bh86_w51_23_c12 & bh86_w51_22_c12 & bh86_w51_21_c12;
   bh86_w51_35_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_c12(0);
   bh86_w52_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_c12(1);
   bh86_w53_28_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid853: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid853_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_copy854_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid853_Out0_copy854_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid855_In0_c12 <= "" & bh86_w51_26_c12 & bh86_w51_27_c12 & bh86_w51_28_c12;
   bh86_w51_36_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_c12(0);
   bh86_w52_32_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid855: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid855_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_copy856_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid855_Out0_copy856_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid857_In0_c12 <= "" & bh86_w52_13_c12 & bh86_w52_28_c12 & bh86_w52_21_c12 & bh86_w52_26_c12 & bh86_w52_20_c12 & bh86_w52_22_c12;
   bh86_w52_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_c12(0);
   bh86_w53_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_c12(1);
   bh86_w54_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid857: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid857_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_copy858_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid857_Out0_copy858_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid859_In0_c12 <= "" & bh86_w52_25_c12 & bh86_w52_27_c12 & bh86_w52_24_c12 & bh86_w52_23_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c0 <= "" & "0";
   bh86_w52_34_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_c12(0);
   bh86_w53_30_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_c12(1);
   bh86_w54_26_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid859: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid859_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid859_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_copy860_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid859_Out0_copy860_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid861_In0_c12 <= "" & bh86_w53_27_c12 & bh86_w53_24_c12 & bh86_w53_25_c12 & bh86_w53_19_c12 & bh86_w53_20_c12 & bh86_w53_21_c12;
   bh86_w53_31_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_c12(0);
   bh86_w54_27_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_c12(1);
   bh86_w55_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid861: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid861_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_copy862_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid861_Out0_copy862_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid863_In0_c12 <= "" & bh86_w53_22_c12 & bh86_w53_23_c12 & bh86_w53_26_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid863_In1_c12 <= "" & bh86_w54_19_c12 & bh86_w54_22_c12;
   bh86_w53_32_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_c12(0);
   bh86_w54_28_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_c12(1);
   bh86_w55_23_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid863: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid863_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid863_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_copy864_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid863_Out0_copy864_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid865_In0_c12 <= "" & bh86_w54_24_c12 & bh86_w54_17_c12 & bh86_w54_18_c12 & bh86_w54_20_c12 & bh86_w54_21_c12 & bh86_w54_23_c12;
   bh86_w54_29_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_c12(0);
   bh86_w55_24_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_c12(1);
   bh86_w56_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid865: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid865_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_copy866_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid865_Out0_copy866_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid867_In0_c12 <= "" & bh86_w55_17_c12 & bh86_w55_21_c12 & bh86_w55_20_c12 & bh86_w55_19_c12 & bh86_w55_18_c12 & bh86_w55_16_c12;
   bh86_w55_25_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_c12(0);
   bh86_w56_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_c12(1);
   bh86_w57_20_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid867: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid867_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_copy868_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid867_Out0_copy868_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid869_In0_c12 <= "" & bh86_w56_20_c12 & bh86_w56_19_c12 & bh86_w56_18_c12 & bh86_w56_17_c12 & bh86_w56_16_c12 & bh86_w56_15_c12;
   bh86_w56_23_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_c12(0);
   bh86_w57_21_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_c12(1);
   bh86_w58_17_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid869: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid869_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_copy870_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid869_Out0_copy870_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid871_In0_c12 <= "" & bh86_w57_19_c12 & bh86_w57_18_c12 & bh86_w57_17_c12 & bh86_w57_16_c12 & bh86_w57_15_c12 & bh86_w57_14_c12;
   bh86_w57_22_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_c12(0);
   bh86_w58_18_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_c12(1);
   bh86_w59_18_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid871: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid871_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_copy872_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid871_Out0_copy872_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid873_In0_c12 <= "" & bh86_w58_11_c12 & bh86_w58_15_c12 & bh86_w58_16_c12 & bh86_w58_14_c12 & bh86_w58_13_c12 & bh86_w58_12_c12;
   bh86_w58_19_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_c12(0);
   bh86_w59_19_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_c12(1);
   bh86_w60_15_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid873: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid873_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_copy874_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid873_Out0_copy874_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid875_In0_c12 <= "" & bh86_w59_17_c12 & bh86_w59_14_c12 & bh86_w59_16_c12 & bh86_w59_15_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid875_In1_c11 <= "" & bh86_w60_10_c11;
   bh86_w59_20_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_c12(0);
   bh86_w60_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_c12(1);
   bh86_w61_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid875: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid875_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid875_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_copy876_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid875_Out0_copy876_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid877_In0_c12 <= "" & bh86_w60_13_c12 & bh86_w60_14_c12 & bh86_w60_12_c12 & bh86_w60_11_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c0 <= "" & "0";
   bh86_w60_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_c12(0);
   bh86_w61_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_c12(1);
   bh86_w62_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid877: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid877_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid877_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_copy878_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid877_Out0_copy878_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid879_In0_c12 <= "" & bh86_w61_12_c12 & bh86_w61_11_c12 & bh86_w61_10_c12;
   bh86_w61_15_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_c12(0);
   bh86_w62_14_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid879: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid879_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_copy880_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid879_Out0_copy880_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid881_In0_c12 <= "" & bh86_w62_12_c12 & bh86_w62_11_c12 & bh86_w62_10_c12;
   bh86_w62_15_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_c12(0);
   bh86_w63_12_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid881: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid881_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_copy882_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid881_Out0_copy882_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid883_In0_c12 <= "" & bh86_w63_8_c12 & bh86_w63_11_c12 & bh86_w63_10_c12 & bh86_w63_9_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c0 <= "" & "0";
   bh86_w63_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_c12(0);
   bh86_w64_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_c12(1);
   bh86_w65_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid883: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid883_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid883_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_copy884_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid883_Out0_copy884_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid885_In0_c12 <= "" & bh86_w64_10_c12 & bh86_w64_9_c12 & bh86_w64_8_c12;
   bh86_w64_12_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_c12(0);
   bh86_w65_13_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid885: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid885_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_copy886_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid885_Out0_copy886_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid887_In0_c12 <= "" & bh86_w65_8_c12 & bh86_w65_11_c12 & bh86_w65_10_c12 & bh86_w65_9_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid887_In1_c12 <= "" & bh86_w66_9_c12;
   bh86_w65_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_c12(0);
   bh86_w66_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_c12(1);
   bh86_w67_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid887: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid887_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid887_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_copy888_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid887_Out0_copy888_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid889_In0_c12 <= "" & bh86_w67_8_c12 & bh86_w67_11_c12 & bh86_w67_10_c12 & bh86_w67_9_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid889_In1_c12 <= "" & bh86_w68_10_c12;
   bh86_w67_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_c12(0);
   bh86_w68_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_c12(1);
   bh86_w69_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid889: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid889_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid889_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_copy890_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid889_Out0_copy890_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid891_In0_c12 <= "" & bh86_w69_10_c12 & bh86_w69_9_c12 & bh86_w69_8_c12;
   bh86_w69_12_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_c12(0);
   bh86_w70_12_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid891: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid891_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_copy892_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid891_Out0_copy892_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid893_In0_c12 <= "" & bh86_w70_8_c12 & bh86_w70_11_c12 & bh86_w70_10_c12 & bh86_w70_9_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid893_In1_c12 <= "" & bh86_w71_9_c12;
   bh86_w70_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_c12(0);
   bh86_w71_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_c12(1);
   bh86_w72_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid893: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid893_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid893_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_copy894_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid893_Out0_copy894_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid895_In0_c12 <= "" & bh86_w72_10_c12 & bh86_w72_9_c12 & bh86_w72_8_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid895_In1_c12 <= "" & bh86_w73_10_c12 & bh86_w73_9_c12;
   bh86_w72_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_c12(0);
   bh86_w73_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_c12(1);
   bh86_w74_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid895: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid895_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid895_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_copy896_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid895_Out0_copy896_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid897_In0_c12 <= "" & bh86_w74_10_c12 & bh86_w74_9_c12 & bh86_w74_8_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c0 <= "" & "0" & "0";
   bh86_w74_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_c12(0);
   bh86_w75_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_c12(1);
   bh86_w76_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid897: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid897_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid897_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_copy898_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid897_Out0_copy898_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid899_In0_c12 <= "" & bh86_w75_10_c12 & bh86_w75_9_c12 & bh86_w75_8_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid899_In1_c12 <= "" & bh86_w76_10_c12 & bh86_w76_9_c12;
   bh86_w75_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_c12(0);
   bh86_w76_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_c12(1);
   bh86_w77_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid899: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid899_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid899_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_copy900_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid899_Out0_copy900_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid901_In0_c12 <= "" & bh86_w77_10_c12 & bh86_w77_9_c12 & bh86_w77_8_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c0 <= "" & "0" & "0";
   bh86_w77_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_c12(0);
   bh86_w78_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_c12(1);
   bh86_w79_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid901: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid901_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid901_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_copy902_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid901_Out0_copy902_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid903_In0_c12 <= "" & bh86_w78_10_c12 & bh86_w78_9_c12 & bh86_w78_8_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid903_In1_c12 <= "" & bh86_w79_10_c12 & bh86_w79_9_c12;
   bh86_w78_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_c12(0);
   bh86_w79_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_c12(1);
   bh86_w80_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid903: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid903_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid903_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_copy904_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid903_Out0_copy904_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid905_In0_c12 <= "" & bh86_w80_10_c12 & bh86_w80_9_c12 & bh86_w80_8_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c0 <= "" & "0" & "0";
   bh86_w80_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_c12(0);
   bh86_w81_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_c12(1);
   bh86_w82_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid905: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid905_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid905_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_copy906_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid905_Out0_copy906_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid907_In0_c12 <= "" & bh86_w81_9_c12 & bh86_w81_8_c12 & bh86_w81_7_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid907_In1_c12 <= "" & bh86_w82_9_c12 & bh86_w82_8_c12;
   bh86_w81_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_c12(0);
   bh86_w82_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_c12(1);
   bh86_w83_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid907: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid907_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid907_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_copy908_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid907_Out0_copy908_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid909_In0_c12 <= "" & bh86_w83_9_c12 & bh86_w83_8_c12 & bh86_w83_7_c12;
   bh86_w83_11_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_c12(0);
   bh86_w84_11_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid909: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid909_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_copy910_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid909_Out0_copy910_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid911_In0_c12 <= "" & bh86_w84_7_c12 & bh86_w84_10_c12 & bh86_w84_9_c12 & bh86_w84_8_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid911_In1_c12 <= "" & bh86_w85_9_c12;
   bh86_w84_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_c12(0);
   bh86_w85_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_c12(1);
   bh86_w86_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid911: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid911_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid911_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_copy912_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid911_Out0_copy912_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid913_In0_c12 <= "" & bh86_w86_9_c12 & bh86_w86_8_c12 & bh86_w86_7_c12;
   bh86_w86_11_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_c12(0);
   bh86_w87_11_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid913: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid913_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_copy914_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid913_Out0_copy914_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid915_In0_c12 <= "" & bh86_w87_7_c12 & bh86_w87_10_c12 & bh86_w87_9_c12 & bh86_w87_8_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid915_In1_c12 <= "" & bh86_w88_8_c12;
   bh86_w87_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_c12(0);
   bh86_w88_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_c12(1);
   bh86_w89_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid915: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid915_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid915_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_copy916_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid915_Out0_copy916_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid917_In0_c12 <= "" & bh86_w89_9_c12 & bh86_w89_8_c12 & bh86_w89_7_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid917_In1_c12 <= "" & bh86_w90_9_c12 & bh86_w90_8_c12;
   bh86_w89_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_c12(0);
   bh86_w90_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_c12(1);
   bh86_w91_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid917: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid917_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid917_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_copy918_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid917_Out0_copy918_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid919_In0_c12 <= "" & bh86_w91_8_c12 & bh86_w91_7_c12 & bh86_w91_6_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c0 <= "" & "0" & "0";
   bh86_w91_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_c12(0);
   bh86_w92_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_c12(1);
   bh86_w93_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid919: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid919_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid919_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_copy920_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid919_Out0_copy920_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid921_In0_c12 <= "" & bh86_w92_8_c12 & bh86_w92_7_c12 & bh86_w92_6_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid921_In1_c12 <= "" & bh86_w93_8_c12 & bh86_w93_7_c12;
   bh86_w92_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_c12(0);
   bh86_w93_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_c12(1);
   bh86_w94_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid921: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid921_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid921_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_copy922_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid921_Out0_copy922_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid923_In0_c12 <= "" & bh86_w94_8_c12 & bh86_w94_7_c12 & bh86_w94_6_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c0 <= "" & "0" & "0";
   bh86_w94_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_c12(0);
   bh86_w95_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_c12(1);
   bh86_w96_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid923: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid923_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid923_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_copy924_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid923_Out0_copy924_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid925_In0_c12 <= "" & bh86_w95_8_c12 & bh86_w95_7_c12 & bh86_w95_6_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid925_In1_c12 <= "" & bh86_w96_8_c12 & bh86_w96_7_c12;
   bh86_w95_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_c12(0);
   bh86_w96_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_c12(1);
   bh86_w97_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid925: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid925_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid925_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_copy926_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid925_Out0_copy926_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid927_In0_c12 <= "" & bh86_w97_8_c12 & bh86_w97_7_c12 & bh86_w97_6_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c0 <= "" & "0" & "0";
   bh86_w97_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_c12(0);
   bh86_w98_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_c12(1);
   bh86_w99_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid927: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid927_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid927_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_copy928_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid927_Out0_copy928_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid929_In0_c12 <= "" & bh86_w98_7_c12 & bh86_w98_6_c12 & bh86_w98_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid929_In1_c12 <= "" & bh86_w99_7_c12 & bh86_w99_6_c12;
   bh86_w98_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_c12(0);
   bh86_w99_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_c12(1);
   bh86_w100_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid929: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid929_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid929_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_copy930_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid929_Out0_copy930_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid931_In0_c12 <= "" & bh86_w100_7_c12 & bh86_w100_6_c12 & bh86_w100_5_c12;
   bh86_w100_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_c12(0);
   bh86_w101_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid931: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid931_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_copy932_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid931_Out0_copy932_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid933_In0_c12 <= "" & bh86_w101_5_c12 & bh86_w101_8_c12 & bh86_w101_7_c12 & bh86_w101_6_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid933_In1_c12 <= "" & bh86_w102_7_c12;
   bh86_w101_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_c12(0);
   bh86_w102_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_c12(1);
   bh86_w103_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid933: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid933_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid933_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_copy934_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid933_Out0_copy934_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid935_In0_c12 <= "" & bh86_w103_7_c12 & bh86_w103_6_c12 & bh86_w103_5_c12;
   bh86_w103_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_c12(0);
   bh86_w104_9_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid935: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid935_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_copy936_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid935_Out0_copy936_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid937_In0_c12 <= "" & bh86_w104_5_c12 & bh86_w104_8_c12 & bh86_w104_7_c12 & bh86_w104_6_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid937_In1_c12 <= "" & bh86_w105_6_c12;
   bh86_w104_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_c12(0);
   bh86_w105_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_c12(1);
   bh86_w106_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid937: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid937_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid937_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_copy938_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid937_Out0_copy938_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid939_In0_c12 <= "" & bh86_w106_7_c12 & bh86_w106_6_c12 & bh86_w106_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid939_In1_c12 <= "" & bh86_w107_7_c12 & bh86_w107_6_c12;
   bh86_w106_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_c12(0);
   bh86_w107_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_c12(1);
   bh86_w108_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid939: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid939_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid939_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_copy940_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid939_Out0_copy940_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid941_In0_c12 <= "" & bh86_w108_7_c12 & bh86_w108_6_c12 & bh86_w108_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c0 <= "" & "0" & "0";
   bh86_w108_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_c12(0);
   bh86_w109_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_c12(1);
   bh86_w110_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid941: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid941_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid941_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_copy942_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid941_Out0_copy942_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid943_In0_c12 <= "" & bh86_w109_7_c12 & bh86_w109_6_c12 & bh86_w109_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid943_In1_c12 <= "" & bh86_w110_7_c12 & bh86_w110_6_c12;
   bh86_w109_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_c12(0);
   bh86_w110_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_c12(1);
   bh86_w111_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid943: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid943_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid943_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_copy944_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid943_Out0_copy944_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid945_In0_c12 <= "" & bh86_w111_7_c12 & bh86_w111_6_c12 & bh86_w111_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c0 <= "" & "0" & "0";
   bh86_w111_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_c12(0);
   bh86_w112_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_c12(1);
   bh86_w113_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid945: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid945_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid945_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_copy946_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid945_Out0_copy946_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid947_In0_c12 <= "" & bh86_w112_7_c12 & bh86_w112_6_c12 & bh86_w112_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid947_In1_c12 <= "" & bh86_w113_7_c12 & bh86_w113_6_c12;
   bh86_w112_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_c12(0);
   bh86_w113_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_c12(1);
   bh86_w114_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid947: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid947_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid947_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_copy948_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid947_Out0_copy948_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid949_In0_c12 <= "" & bh86_w114_7_c12 & bh86_w114_6_c12 & bh86_w114_5_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid949_In1_c12 <= "" & bh86_w115_2_c12 & bh86_w115_4_c12;
   bh86_w114_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_c12(0);
   bh86_w115_5_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_c12(1);
   bh86_w116_5_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid949: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid949_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid949_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_copy950_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid949_Out0_copy950_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid951_In0_c12 <= "" & bh86_w116_4_c12 & bh86_w116_3_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid951_In1_c12 <= "" & bh86_w117_2_c12;
   bh86_w116_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_c12(0);
   bh86_w117_3_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_c12(1);
   bh86_w118_2_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid951: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid951_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid951_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_copy952_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid951_Out0_copy952_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid953_In0_c12 <= "" & bh86_w118_0_c12 & bh86_w118_1_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid953_In1_c11 <= "" & bh86_w119_0_c11;
   bh86_w118_3_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_c12(0);
   bh86_w119_1_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_c12(1);
   Compressor_14_3_Freq300_uid626_uid953: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid953_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid953_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_copy954_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid953_Out0_copy954_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid955_In0_c12 <= "" & bh86_w45_29_c12 & bh86_w45_30_c12 & bh86_w45_31_c12;
   bh86_w45_32_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_c12(0);
   bh86_w46_37_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid955: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid955_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_copy956_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid955_Out0_copy956_c12; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid959_In0_c12 <= "" & bh86_w46_33_c12 & bh86_w46_35_c12 & bh86_w46_32_c12 & bh86_w46_34_c12 & bh86_w46_36_c12;
   bh86_w46_38_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_c12(0);
   bh86_w47_41_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_c12(1);
   bh86_w48_40_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_c12(2);
   Compressor_5_3_Freq300_uid958_uid959: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid959_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_copy960_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid959_Out0_copy960_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid961_In0_c12 <= "" & bh86_w47_40_c12 & bh86_w47_36_c12 & bh86_w47_37_c12 & bh86_w47_39_c12 & bh86_w47_26_c12 & bh86_w47_38_c12;
   bh86_w47_42_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_c12(0);
   bh86_w48_41_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_c12(1);
   bh86_w49_41_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid961: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid961_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_copy962_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid961_Out0_copy962_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid963_In0_c12 <= "" & bh86_w48_36_c12 & bh86_w48_37_c12 & bh86_w48_34_c12 & bh86_w48_23_c12 & bh86_w48_39_c12 & bh86_w48_38_c12;
   bh86_w48_42_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_c12(0);
   bh86_w49_42_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_c12(1);
   bh86_w50_38_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid963: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid963_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_copy964_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid963_Out0_copy964_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid965_In0_c12 <= "" & bh86_w49_39_c12 & bh86_w49_36_c12 & bh86_w49_35_c12 & bh86_w49_38_c12 & bh86_w49_40_c12 & bh86_w49_37_c12;
   bh86_w49_43_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_c12(0);
   bh86_w50_39_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_c12(1);
   bh86_w51_37_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid965: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid965_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_copy966_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid965_Out0_copy966_c12; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid967_In0_c12 <= "" & bh86_w50_34_c12 & bh86_w50_37_c12 & bh86_w50_36_c12 & bh86_w50_33_c12 & bh86_w50_35_c12;
   bh86_w50_40_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_c12(0);
   bh86_w51_38_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_c12(1);
   bh86_w52_35_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_c12(2);
   Compressor_5_3_Freq300_uid958_uid967: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid967_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_copy968_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_c12 <= Compressor_5_3_Freq300_uid958_bh86_uid967_Out0_copy968_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid969_In0_c12 <= "" & bh86_w51_31_c12 & bh86_w51_36_c12 & bh86_w51_34_c12 & bh86_w51_35_c12 & bh86_w51_32_c12 & bh86_w51_33_c12;
   bh86_w51_39_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_c12(0);
   bh86_w52_36_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_c12(1);
   bh86_w53_33_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid969: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid969_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_copy970_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid969_Out0_copy970_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid971_In0_c12 <= "" & bh86_w52_34_c12 & bh86_w52_32_c12 & bh86_w52_30_c12 & bh86_w52_33_c12 & bh86_w52_31_c12 & bh86_w52_29_c12;
   bh86_w52_37_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_c12(0);
   bh86_w53_34_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_c12(1);
   bh86_w54_30_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_c12(2);
   Compressor_6_3_Freq300_uid616_uid971: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid971_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_copy972_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_c12 <= Compressor_6_3_Freq300_uid616_bh86_uid971_Out0_copy972_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid973_In0_c12 <= "" & bh86_w53_30_c12 & bh86_w53_32_c12 & bh86_w53_31_c12 & bh86_w53_29_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid973_In1_c12 <= "" & bh86_w54_26_c12;
   bh86_w53_35_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_c12(0);
   bh86_w54_31_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_c12(1);
   bh86_w55_26_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid973: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid973_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid973_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_copy974_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid973_Out0_copy974_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid975_In0_c12 <= "" & bh86_w54_28_c12 & bh86_w54_29_c12 & bh86_w54_27_c12 & bh86_w54_25_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid975_In1_c12 <= "" & bh86_w55_15_c12;
   bh86_w54_32_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_c12(0);
   bh86_w55_27_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_c12(1);
   bh86_w56_24_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid975: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid975_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid975_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_copy976_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid975_Out0_copy976_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid977_In0_c12 <= "" & bh86_w55_23_c12 & bh86_w55_25_c12 & bh86_w55_24_c12 & bh86_w55_22_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c0 <= "" & "0";
   bh86_w55_28_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_c12(0);
   bh86_w56_25_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_c12(1);
   bh86_w57_23_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid977: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid977_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid977_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_copy978_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid977_Out0_copy978_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid979_In0_c12 <= "" & bh86_w56_23_c12 & bh86_w56_22_c12 & bh86_w56_21_c12;
   bh86_w56_26_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_c12(0);
   bh86_w57_24_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid979: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid979_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_copy980_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid979_Out0_copy980_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid981_In0_c12 <= "" & bh86_w57_22_c12 & bh86_w57_21_c12 & bh86_w57_20_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid981_In1_c12 <= "" & bh86_w58_19_c12 & bh86_w58_18_c12;
   bh86_w57_25_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_c12(0);
   bh86_w58_20_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_c12(1);
   bh86_w59_21_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid981: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid981_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid981_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_copy982_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid981_Out0_copy982_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid983_In0_c12 <= "" & bh86_w59_13_c12 & bh86_w59_20_c12 & bh86_w59_19_c12 & bh86_w59_18_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c0 <= "" & "0";
   bh86_w59_22_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_c12(0);
   bh86_w60_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_c12(1);
   bh86_w61_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid983: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid983_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid983_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_copy984_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid983_Out0_copy984_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid985_In0_c12 <= "" & bh86_w60_17_c12 & bh86_w60_16_c12 & bh86_w60_15_c12;
   bh86_w60_19_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_c12(0);
   bh86_w61_17_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid985: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid985_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_copy986_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid985_Out0_copy986_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid987_In0_c12 <= "" & bh86_w61_14_c12 & bh86_w61_15_c12 & bh86_w61_13_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid987_In1_c12 <= "" & bh86_w62_13_c12 & bh86_w62_15_c12;
   bh86_w61_18_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_c12(0);
   bh86_w62_16_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_c12(1);
   bh86_w63_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid987: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid987_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid987_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_copy988_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid987_Out0_copy988_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid989_In0_c12 <= "" & bh86_w63_13_c12 & bh86_w63_12_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid989_In1_c12 <= "" & bh86_w64_11_c12 & bh86_w64_12_c12;
   bh86_w63_15_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_c12(0);
   bh86_w64_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_c12(1);
   bh86_w65_15_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid989: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid989_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid989_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_copy990_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid989_Out0_copy990_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid991_In0_c12 <= "" & bh86_w65_12_c12 & bh86_w65_14_c12 & bh86_w65_13_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid991_In1_c12 <= "" & bh86_w66_8_c12 & bh86_w66_10_c12;
   bh86_w65_16_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_c12(0);
   bh86_w66_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_c12(1);
   bh86_w67_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid991: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid991_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid991_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_copy992_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid991_Out0_copy992_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid993_In0_c12 <= "" & bh86_w67_13_c12 & bh86_w67_12_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid993_In1_c12 <= "" & bh86_w68_9_c12 & bh86_w68_11_c12;
   bh86_w67_15_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_c12(0);
   bh86_w68_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_c12(1);
   bh86_w69_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid993: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid993_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid993_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_copy994_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid993_Out0_copy994_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid995_In0_c12 <= "" & bh86_w69_12_c12 & bh86_w69_11_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid995_In1_c12 <= "" & bh86_w70_13_c12 & bh86_w70_12_c12;
   bh86_w69_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_c12(0);
   bh86_w70_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_c12(1);
   bh86_w71_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid995: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid995_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid995_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_copy996_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid995_Out0_copy996_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid997_In0_c12 <= "" & bh86_w71_8_c12 & bh86_w71_10_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid997_In1_c12 <= "" & bh86_w72_12_c12 & bh86_w72_11_c12;
   bh86_w71_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_c12(0);
   bh86_w72_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_c12(1);
   bh86_w73_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid997: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid997_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid997_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_copy998_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid997_Out0_copy998_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid999_In0_c12 <= "" & bh86_w74_12_c12 & bh86_w74_11_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid999_In1_c12 <= "" & bh86_w75_11_c12 & bh86_w75_12_c12;
   bh86_w74_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_c12(0);
   bh86_w75_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_c12(1);
   bh86_w76_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid999: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid999_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid999_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_copy1000_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid999_Out0_copy1000_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1001_In0_c12 <= "" & bh86_w76_11_c12 & bh86_w76_12_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1001_In1_c12 <= "" & bh86_w77_12_c12 & bh86_w77_11_c12;
   bh86_w76_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_c12(0);
   bh86_w77_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_c12(1);
   bh86_w78_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1001: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1001_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1001_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_copy1002_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1001_Out0_copy1002_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1003_In0_c12 <= "" & bh86_w78_11_c12 & bh86_w78_12_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1003_In1_c12 <= "" & bh86_w79_11_c12 & bh86_w79_12_c12;
   bh86_w78_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_c12(0);
   bh86_w79_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_c12(1);
   bh86_w80_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1003: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1003_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1003_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_copy1004_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1003_Out0_copy1004_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1005_In0_c12 <= "" & bh86_w80_12_c12 & bh86_w80_11_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1005_In1_c12 <= "" & bh86_w81_10_c12 & bh86_w81_11_c12;
   bh86_w80_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_c12(0);
   bh86_w81_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_c12(1);
   bh86_w82_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1005: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1005_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1005_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_copy1006_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1005_Out0_copy1006_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1007_In0_c12 <= "" & bh86_w82_10_c12 & bh86_w82_11_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1007_In1_c12 <= "" & bh86_w83_11_c12 & bh86_w83_10_c12;
   bh86_w82_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_c12(0);
   bh86_w83_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_c12(1);
   bh86_w84_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1007: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1007_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1007_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_copy1008_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1007_Out0_copy1008_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1009_In0_c12 <= "" & bh86_w84_12_c12 & bh86_w84_11_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1009_In1_c12 <= "" & bh86_w85_8_c12 & bh86_w85_10_c12;
   bh86_w84_14_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_c12(0);
   bh86_w85_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_c12(1);
   bh86_w86_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1009: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1009_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1009_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_copy1010_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1009_Out0_copy1010_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1011_In0_c12 <= "" & bh86_w86_11_c12 & bh86_w86_10_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1011_In1_c12 <= "" & bh86_w87_12_c12 & bh86_w87_11_c12;
   bh86_w86_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_c12(0);
   bh86_w87_13_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_c12(1);
   bh86_w88_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1011: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1011_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1011_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_copy1012_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1011_Out0_copy1012_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1013_In0_c12 <= "" & bh86_w88_7_c12 & bh86_w88_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1013_In1_c12 <= "" & bh86_w89_11_c12 & bh86_w89_10_c12;
   bh86_w88_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_c12(0);
   bh86_w89_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_c12(1);
   bh86_w90_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1013: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1013_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1013_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_copy1014_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1013_Out0_copy1014_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1015_In0_c12 <= "" & bh86_w91_10_c12 & bh86_w91_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1015_In1_c12 <= "" & bh86_w92_9_c12 & bh86_w92_10_c12;
   bh86_w91_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_c12(0);
   bh86_w92_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_c12(1);
   bh86_w93_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1015: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1015_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1015_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_copy1016_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1015_Out0_copy1016_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1017_In0_c12 <= "" & bh86_w93_9_c12 & bh86_w93_10_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1017_In1_c12 <= "" & bh86_w94_10_c12 & bh86_w94_9_c12;
   bh86_w93_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_c12(0);
   bh86_w94_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_c12(1);
   bh86_w95_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1017: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1017_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1017_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_copy1018_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1017_Out0_copy1018_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1019_In0_c12 <= "" & bh86_w95_9_c12 & bh86_w95_10_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1019_In1_c12 <= "" & bh86_w96_9_c12 & bh86_w96_10_c12;
   bh86_w95_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_c12(0);
   bh86_w96_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_c12(1);
   bh86_w97_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1019: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1019_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1019_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_copy1020_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1019_Out0_copy1020_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1021_In0_c12 <= "" & bh86_w97_10_c12 & bh86_w97_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1021_In1_c12 <= "" & bh86_w98_8_c12 & bh86_w98_9_c12;
   bh86_w97_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_c12(0);
   bh86_w98_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_c12(1);
   bh86_w99_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1021: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1021_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1021_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_copy1022_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1021_Out0_copy1022_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1023_In0_c12 <= "" & bh86_w99_8_c12 & bh86_w99_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1023_In1_c12 <= "" & bh86_w100_9_c12 & bh86_w100_8_c12;
   bh86_w99_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_c12(0);
   bh86_w100_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_c12(1);
   bh86_w101_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1023: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1023_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1023_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_copy1024_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1023_Out0_copy1024_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1025_In0_c12 <= "" & bh86_w101_10_c12 & bh86_w101_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1025_In1_c12 <= "" & bh86_w102_6_c12 & bh86_w102_8_c12;
   bh86_w101_12_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_c12(0);
   bh86_w102_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_c12(1);
   bh86_w103_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1025: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1025_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1025_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_copy1026_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1025_Out0_copy1026_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1027_In0_c12 <= "" & bh86_w103_9_c12 & bh86_w103_8_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1027_In1_c12 <= "" & bh86_w104_10_c12 & bh86_w104_9_c12;
   bh86_w103_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_c12(0);
   bh86_w104_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_c12(1);
   bh86_w105_8_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1027: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1027_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1027_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_copy1028_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1027_Out0_copy1028_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1029_In0_c12 <= "" & bh86_w105_5_c12 & bh86_w105_7_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1029_In1_c12 <= "" & bh86_w106_9_c12 & bh86_w106_8_c12;
   bh86_w105_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_c12(0);
   bh86_w106_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_c12(1);
   bh86_w107_9_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1029: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1029_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1029_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_copy1030_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1029_Out0_copy1030_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1031_In0_c12 <= "" & bh86_w108_9_c12 & bh86_w108_8_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1031_In1_c12 <= "" & bh86_w109_8_c12 & bh86_w109_9_c12;
   bh86_w108_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_c12(0);
   bh86_w109_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_c12(1);
   bh86_w110_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1031: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1031_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1031_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_copy1032_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1031_Out0_copy1032_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1033_In0_c12 <= "" & bh86_w110_8_c12 & bh86_w110_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1033_In1_c12 <= "" & bh86_w111_9_c12 & bh86_w111_8_c12;
   bh86_w110_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_c12(0);
   bh86_w111_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_c12(1);
   bh86_w112_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1033: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1033_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1033_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_copy1034_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1033_Out0_copy1034_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1035_In0_c12 <= "" & bh86_w112_8_c12 & bh86_w112_9_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1035_In1_c12 <= "" & bh86_w113_8_c12 & bh86_w113_9_c12;
   bh86_w112_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_c12(0);
   bh86_w113_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_c12(1);
   bh86_w114_10_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1035: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1035_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1035_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_copy1036_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1035_Out0_copy1036_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1037_In0_c12 <= "" & bh86_w114_9_c12 & bh86_w114_8_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1037_In1_c12 <= "" & bh86_w115_3_c12 & bh86_w115_5_c12;
   bh86_w114_11_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_c12(0);
   bh86_w115_6_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_c12(1);
   bh86_w116_7_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1037: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1037_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1037_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_copy1038_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1037_Out0_copy1038_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1039_In0_c12 <= "" & bh86_w116_6_c12 & bh86_w116_5_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1039_In1_c12 <= "" & bh86_w117_3_c12;
   bh86_w116_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_c12(0);
   bh86_w117_4_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_c12(1);
   bh86_w118_4_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1039: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1039_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1039_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_copy1040_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1039_Out0_copy1040_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1041_In0_c12 <= "" & bh86_w118_3_c12 & bh86_w118_2_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1041_In1_c12 <= "" & bh86_w119_1_c12;
   bh86_w118_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_c12(0);
   bh86_w119_2_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_c12(1);
   Compressor_14_3_Freq300_uid626_uid1041: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1041_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1041_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_copy1042_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1041_Out0_copy1042_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1043_In0_c12 <= "" & bh86_w46_37_c12 & bh86_w46_38_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1043_In1_c12 <= "" & bh86_w47_41_c12 & bh86_w47_42_c12;
   bh86_w46_39_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_c12(0);
   bh86_w47_43_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_c12(1);
   bh86_w48_43_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1043: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1043_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1043_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_copy1044_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1043_Out0_copy1044_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1045_In0_c12 <= "" & bh86_w48_40_c12 & bh86_w48_41_c12 & bh86_w48_42_c12 & bh86_w48_35_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c0 <= "" & "0";
   bh86_w48_44_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_c12(0);
   bh86_w49_44_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_c12(1);
   bh86_w50_41_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1045: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1045_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1045_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_copy1046_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1045_Out0_copy1046_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1047_In0_c12 <= "" & bh86_w49_41_c12 & bh86_w49_42_c12 & bh86_w49_43_c12;
   bh86_w49_45_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_c12(0);
   bh86_w50_42_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1047: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1047_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_copy1048_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1047_Out0_copy1048_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1049_In0_c12 <= "" & bh86_w50_38_c12 & bh86_w50_39_c12 & bh86_w50_40_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1049_In1_c12 <= "" & bh86_w51_37_c12 & bh86_w51_38_c12;
   bh86_w50_43_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_c12(0);
   bh86_w51_40_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_c12(1);
   bh86_w52_38_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1049: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1049_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1049_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_copy1050_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1049_Out0_copy1050_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1051_In0_c12 <= "" & bh86_w52_35_c12 & bh86_w52_36_c12 & bh86_w52_37_c12;
   bh86_w52_39_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_c12(0);
   bh86_w53_36_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1051: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1051_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_copy1052_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1051_Out0_copy1052_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1053_In0_c12 <= "" & bh86_w53_33_c12 & bh86_w53_34_c12 & bh86_w53_35_c12 & bh86_w53_28_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c0 <= "" & "0";
   bh86_w53_37_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_c12(0);
   bh86_w54_33_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_c12(1);
   bh86_w55_29_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1053: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1053_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1053_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_copy1054_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1053_Out0_copy1054_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1055_In0_c12 <= "" & bh86_w54_30_c12 & bh86_w54_31_c12 & bh86_w54_32_c12;
   bh86_w54_34_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_c12(0);
   bh86_w55_30_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1055: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1055_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_copy1056_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1055_Out0_copy1056_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1057_In0_c12 <= "" & bh86_w55_26_c12 & bh86_w55_28_c12 & bh86_w55_27_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1057_In1_c12 <= "" & bh86_w56_25_c12 & bh86_w56_26_c12;
   bh86_w55_31_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_c12(0);
   bh86_w56_27_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_c12(1);
   bh86_w57_26_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1057: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1057_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1057_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_copy1058_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1057_Out0_copy1058_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1059_In0_c12 <= "" & bh86_w57_23_c12 & bh86_w57_25_c12 & bh86_w57_24_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1059_In1_c12 <= "" & bh86_w58_17_c12 & bh86_w58_20_c12;
   bh86_w57_27_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_c12(0);
   bh86_w58_21_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_c12(1);
   bh86_w59_23_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1059: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1059_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1059_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_copy1060_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1059_Out0_copy1060_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1061_In0_c12 <= "" & bh86_w59_22_c12 & bh86_w59_21_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1061_In1_c12 <= "" & bh86_w60_18_c12 & bh86_w60_19_c12;
   bh86_w59_24_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_c12(0);
   bh86_w60_20_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_c12(1);
   bh86_w61_19_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1061: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1061_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1061_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_copy1062_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1061_Out0_copy1062_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1063_In0_c12 <= "" & bh86_w61_16_c12 & bh86_w61_17_c12 & bh86_w61_18_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1063_In1_c12 <= "" & bh86_w62_16_c12 & bh86_w62_14_c12;
   bh86_w61_20_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_c12(0);
   bh86_w62_17_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_c12(1);
   bh86_w63_16_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1063: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1063_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1063_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_copy1064_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1063_Out0_copy1064_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1065_In0_c12 <= "" & bh86_w63_14_c12 & bh86_w63_15_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1065_In1_c12 <= "" & bh86_w64_13_c12;
   bh86_w63_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_c12(0);
   bh86_w64_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_c12(1);
   bh86_w65_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1065: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1065_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1065_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_copy1066_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1065_Out0_copy1066_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1067_In0_c12 <= "" & bh86_w65_15_c12 & bh86_w65_16_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1067_In1_c12 <= "" & bh86_w66_11_c12;
   bh86_w65_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_c12(0);
   bh86_w66_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_c12(1);
   bh86_w67_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1067: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1067_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1067_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_copy1068_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1067_Out0_copy1068_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1069_In0_c12 <= "" & bh86_w67_14_c12 & bh86_w67_15_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1069_In1_c12 <= "" & bh86_w68_12_c12;
   bh86_w67_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_c12(0);
   bh86_w68_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_c12(1);
   bh86_w69_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1069: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1069_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1069_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_copy1070_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1069_Out0_copy1070_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1071_In0_c12 <= "" & bh86_w69_14_c12 & bh86_w69_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1071_In1_c12 <= "" & bh86_w70_14_c12;
   bh86_w69_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_c12(0);
   bh86_w70_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_c12(1);
   bh86_w71_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1071: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1071_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1071_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_copy1072_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1071_Out0_copy1072_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1073_In0_c12 <= "" & bh86_w71_12_c12 & bh86_w71_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1073_In1_c12 <= "" & bh86_w72_13_c12;
   bh86_w71_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_c12(0);
   bh86_w72_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_c12(1);
   bh86_w73_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1073: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1073_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1073_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_copy1074_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1073_Out0_copy1074_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1075_In0_c12 <= "" & bh86_w73_11_c12 & bh86_w73_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1075_In1_c12 <= "" & bh86_w74_13_c12;
   bh86_w73_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_c12(0);
   bh86_w74_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_c12(1);
   bh86_w75_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1075: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1075_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1075_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_copy1076_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1075_Out0_copy1076_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1077_In0_c12 <= "" & bh86_w76_13_c12 & bh86_w76_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1077_In1_c12 <= "" & bh86_w77_13_c12;
   bh86_w76_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_c12(0);
   bh86_w77_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_c12(1);
   bh86_w78_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1077: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1077_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1077_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_copy1078_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1077_Out0_copy1078_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1079_In0_c12 <= "" & bh86_w78_13_c12 & bh86_w78_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1079_In1_c12 <= "" & bh86_w79_13_c12;
   bh86_w78_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_c12(0);
   bh86_w79_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_c12(1);
   bh86_w80_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1079: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1079_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1079_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_copy1080_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1079_Out0_copy1080_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1081_In0_c12 <= "" & bh86_w80_13_c12 & bh86_w80_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1081_In1_c12 <= "" & bh86_w81_12_c12;
   bh86_w80_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_c12(0);
   bh86_w81_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_c12(1);
   bh86_w82_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1081: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1081_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1081_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_copy1082_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1081_Out0_copy1082_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1083_In0_c12 <= "" & bh86_w82_12_c12 & bh86_w82_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1083_In1_c12 <= "" & bh86_w83_12_c12;
   bh86_w82_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_c12(0);
   bh86_w83_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_c12(1);
   bh86_w84_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1083: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1083_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1083_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_copy1084_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1083_Out0_copy1084_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1085_In0_c12 <= "" & bh86_w84_13_c12 & bh86_w84_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1085_In1_c12 <= "" & bh86_w85_11_c12;
   bh86_w84_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_c12(0);
   bh86_w85_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_c12(1);
   bh86_w86_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1085: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1085_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1085_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_copy1086_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1085_Out0_copy1086_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1087_In0_c12 <= "" & bh86_w86_13_c12 & bh86_w86_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1087_In1_c12 <= "" & bh86_w87_13_c12;
   bh86_w86_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_c12(0);
   bh86_w87_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_c12(1);
   bh86_w88_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1087: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1087_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1087_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_copy1088_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1087_Out0_copy1088_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1089_In0_c12 <= "" & bh86_w88_11_c12 & bh86_w88_10_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1089_In1_c12 <= "" & bh86_w89_12_c12;
   bh86_w88_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_c12(0);
   bh86_w89_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_c12(1);
   bh86_w90_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1089: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1089_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1089_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_copy1090_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1089_Out0_copy1090_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1091_In0_c12 <= "" & bh86_w90_10_c12 & bh86_w90_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1091_In1_c12 <= "" & bh86_w91_11_c12;
   bh86_w90_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_c12(0);
   bh86_w91_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_c12(1);
   bh86_w92_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1091: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1091_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1091_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_copy1092_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1091_Out0_copy1092_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1093_In0_c12 <= "" & bh86_w93_11_c12 & bh86_w93_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1093_In1_c12 <= "" & bh86_w94_11_c12;
   bh86_w93_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_c12(0);
   bh86_w94_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_c12(1);
   bh86_w95_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1093: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1093_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1093_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_copy1094_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1093_Out0_copy1094_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1095_In0_c12 <= "" & bh86_w95_11_c12 & bh86_w95_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1095_In1_c12 <= "" & bh86_w96_11_c12;
   bh86_w95_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_c12(0);
   bh86_w96_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_c12(1);
   bh86_w97_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1095: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1095_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1095_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_copy1096_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1095_Out0_copy1096_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1097_In0_c12 <= "" & bh86_w97_11_c12 & bh86_w97_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1097_In1_c12 <= "" & bh86_w98_10_c12;
   bh86_w97_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_c12(0);
   bh86_w98_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_c12(1);
   bh86_w99_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1097: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1097_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1097_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_copy1098_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1097_Out0_copy1098_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1099_In0_c12 <= "" & bh86_w99_10_c12 & bh86_w99_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1099_In1_c12 <= "" & bh86_w100_10_c12;
   bh86_w99_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_c12(0);
   bh86_w100_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_c12(1);
   bh86_w101_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1099: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1099_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1099_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_copy1100_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1099_Out0_copy1100_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1101_In0_c12 <= "" & bh86_w101_11_c12 & bh86_w101_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1101_In1_c12 <= "" & bh86_w102_9_c12;
   bh86_w101_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_c12(0);
   bh86_w102_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_c12(1);
   bh86_w103_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1101: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1101_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1101_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_copy1102_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1101_Out0_copy1102_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1103_In0_c12 <= "" & bh86_w103_11_c12 & bh86_w103_10_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1103_In1_c12 <= "" & bh86_w104_11_c12;
   bh86_w103_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_c12(0);
   bh86_w104_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_c12(1);
   bh86_w105_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1103: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1103_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1103_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_copy1104_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1103_Out0_copy1104_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1105_In0_c12 <= "" & bh86_w105_9_c12 & bh86_w105_8_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1105_In1_c12 <= "" & bh86_w106_10_c12;
   bh86_w105_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_c12(0);
   bh86_w106_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_c12(1);
   bh86_w107_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1105: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1105_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1105_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_copy1106_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1105_Out0_copy1106_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1107_In0_c12 <= "" & bh86_w107_8_c12 & bh86_w107_9_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1107_In1_c12 <= "" & bh86_w108_10_c12;
   bh86_w107_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_c12(0);
   bh86_w108_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_c12(1);
   bh86_w109_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1107: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1107_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1107_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_copy1108_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1107_Out0_copy1108_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1109_In0_c12 <= "" & bh86_w110_10_c12 & bh86_w110_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1109_In1_c12 <= "" & bh86_w111_10_c12;
   bh86_w110_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_c12(0);
   bh86_w111_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_c12(1);
   bh86_w112_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1109: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1109_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1109_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_copy1110_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1109_Out0_copy1110_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1111_In0_c12 <= "" & bh86_w112_10_c12 & bh86_w112_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1111_In1_c12 <= "" & bh86_w113_10_c12;
   bh86_w112_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_c12(0);
   bh86_w113_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_c12(1);
   bh86_w114_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1111: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1111_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1111_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_copy1112_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1111_Out0_copy1112_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1113_In0_c12 <= "" & bh86_w114_10_c12 & bh86_w114_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1113_In1_c12 <= "" & bh86_w115_6_c12;
   bh86_w114_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_c12(0);
   bh86_w115_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_c12(1);
   bh86_w116_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1113: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1113_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1113_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_copy1114_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1113_Out0_copy1114_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1115_In0_c12 <= "" & bh86_w116_8_c12 & bh86_w116_7_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1115_In1_c12 <= "" & bh86_w117_4_c12;
   bh86_w116_10_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_c12(0);
   bh86_w117_5_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_c12(1);
   bh86_w118_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1115: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1115_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1115_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_copy1116_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1115_Out0_copy1116_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1117_In0_c12 <= "" & bh86_w118_5_c12 & bh86_w118_4_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1117_In1_c12 <= "" & bh86_w119_2_c12;
   bh86_w118_7_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_c12(0);
   bh86_w119_3_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_c12(1);
   Compressor_14_3_Freq300_uid626_uid1117: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1117_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1117_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_copy1118_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1117_Out0_copy1118_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1119_In0_c12 <= "" & bh86_w48_43_c12 & bh86_w48_44_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1119_In1_c12 <= "" & bh86_w49_44_c12 & bh86_w49_45_c12;
   bh86_w48_45_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_c12(0);
   bh86_w49_46_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_c12(1);
   bh86_w50_44_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1119: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1119_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1119_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_copy1120_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1119_Out0_copy1120_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1121_In0_c12 <= "" & bh86_w50_41_c12 & bh86_w50_42_c12 & bh86_w50_43_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1121_In1_c12 <= "" & bh86_w51_39_c12 & bh86_w51_40_c12;
   bh86_w50_45_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_c12(0);
   bh86_w51_41_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_c12(1);
   bh86_w52_40_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1121: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1121_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1121_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_copy1122_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1121_Out0_copy1122_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1123_In0_c12 <= "" & bh86_w52_38_c12 & bh86_w52_39_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1123_In1_c12 <= "" & bh86_w53_36_c12 & bh86_w53_37_c12;
   bh86_w52_41_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_c12(0);
   bh86_w53_38_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_c12(1);
   bh86_w54_35_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1123: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1123_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1123_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_copy1124_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1123_Out0_copy1124_c12; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1125_In0_c12 <= "" & bh86_w54_33_c12 & bh86_w54_34_c12 & "0";
   bh86_w54_36_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_c12(0);
   bh86_w55_32_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1125: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1125_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_copy1126_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1125_Out0_copy1126_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1127_In0_c12 <= "" & bh86_w55_29_c12 & bh86_w55_30_c12 & bh86_w55_31_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1127_In1_c12 <= "" & bh86_w56_27_c12 & bh86_w56_24_c12;
   bh86_w55_33_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_c12(0);
   bh86_w56_28_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_c12(1);
   bh86_w57_28_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1127: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1127_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1127_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_copy1128_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1127_Out0_copy1128_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1129_In0_c12 <= "" & bh86_w57_26_c12 & bh86_w57_27_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1129_In1_c12 <= "" & bh86_w58_21_c12;
   bh86_w57_29_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_c12(0);
   bh86_w58_22_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_c12(1);
   bh86_w59_25_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1129: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1129_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1129_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_copy1130_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1129_Out0_copy1130_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1131_In0_c12 <= "" & bh86_w59_23_c12 & bh86_w59_24_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1131_In1_c12 <= "" & bh86_w60_20_c12;
   bh86_w59_26_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_c12(0);
   bh86_w60_21_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_c12(1);
   bh86_w61_21_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1131: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1131_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1131_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_copy1132_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1131_Out0_copy1132_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1133_In0_c12 <= "" & bh86_w61_19_c12 & bh86_w61_20_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1133_In1_c12 <= "" & bh86_w62_17_c12;
   bh86_w61_22_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_c12(0);
   bh86_w62_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_c12(1);
   bh86_w63_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1133: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1133_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1133_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_copy1134_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1133_Out0_copy1134_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1135_In0_c12 <= "" & bh86_w63_16_c12 & bh86_w63_17_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1135_In1_c12 <= "" & bh86_w64_14_c12;
   bh86_w63_19_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_c12(0);
   bh86_w64_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_c12(1);
   bh86_w65_19_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1135: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1135_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1135_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_copy1136_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1135_Out0_copy1136_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1137_In0_c12 <= "" & bh86_w65_17_c12 & bh86_w65_18_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1137_In1_c12 <= "" & bh86_w66_12_c12;
   bh86_w65_20_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_c12(0);
   bh86_w66_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_c12(1);
   bh86_w67_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1137: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1137_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1137_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_copy1138_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1137_Out0_copy1138_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1139_In0_c12 <= "" & bh86_w67_16_c12 & bh86_w67_17_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1139_In1_c12 <= "" & bh86_w68_13_c12;
   bh86_w67_19_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_c12(0);
   bh86_w68_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_c12(1);
   bh86_w69_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1139: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1139_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1139_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_copy1140_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1139_Out0_copy1140_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1141_In0_c12 <= "" & bh86_w69_15_c12 & bh86_w69_16_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1141_In1_c12 <= "" & bh86_w70_15_c12;
   bh86_w69_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_c12(0);
   bh86_w70_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_c12(1);
   bh86_w71_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1141: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1141_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1141_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_copy1142_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1141_Out0_copy1142_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1143_In0_c12 <= "" & bh86_w71_14_c12 & bh86_w71_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1143_In1_c12 <= "" & bh86_w72_14_c12;
   bh86_w71_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_c12(0);
   bh86_w72_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_c12(1);
   bh86_w73_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1143: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1143_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1143_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_copy1144_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1143_Out0_copy1144_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1145_In0_c12 <= "" & bh86_w73_14_c12 & bh86_w73_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1145_In1_c12 <= "" & bh86_w74_14_c12;
   bh86_w73_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_c12(0);
   bh86_w74_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_c12(1);
   bh86_w75_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1145: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1145_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1145_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_copy1146_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1145_Out0_copy1146_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1147_In0_c12 <= "" & bh86_w75_13_c12 & bh86_w75_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1147_In1_c12 <= "" & bh86_w76_15_c12;
   bh86_w75_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_c12(0);
   bh86_w76_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_c12(1);
   bh86_w77_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1147: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1147_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1147_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_copy1148_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1147_Out0_copy1148_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1149_In0_c12 <= "" & bh86_w78_15_c12 & bh86_w78_16_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1149_In1_c12 <= "" & bh86_w79_14_c12;
   bh86_w78_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_c12(0);
   bh86_w79_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_c12(1);
   bh86_w80_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1149: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1149_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1149_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_copy1150_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1149_Out0_copy1150_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1151_In0_c12 <= "" & bh86_w80_15_c12 & bh86_w80_16_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1151_In1_c12 <= "" & bh86_w81_13_c12;
   bh86_w80_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_c12(0);
   bh86_w81_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_c12(1);
   bh86_w82_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1151: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1151_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1151_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_copy1152_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1151_Out0_copy1152_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1153_In0_c12 <= "" & bh86_w82_14_c12 & bh86_w82_15_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1153_In1_c12 <= "" & bh86_w83_13_c12;
   bh86_w82_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_c12(0);
   bh86_w83_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_c12(1);
   bh86_w84_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1153: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1153_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1153_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_copy1154_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1153_Out0_copy1154_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1155_In0_c12 <= "" & bh86_w84_15_c12 & bh86_w84_16_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1155_In1_c12 <= "" & bh86_w85_12_c12;
   bh86_w84_18_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_c12(0);
   bh86_w85_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_c12(1);
   bh86_w86_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1155: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1155_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1155_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_copy1156_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1155_Out0_copy1156_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1157_In0_c12 <= "" & bh86_w86_14_c12 & bh86_w86_15_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1157_In1_c12 <= "" & bh86_w87_14_c12;
   bh86_w86_17_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_c12(0);
   bh86_w87_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_c12(1);
   bh86_w88_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1157: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1157_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1157_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_copy1158_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1157_Out0_copy1158_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1159_In0_c12 <= "" & bh86_w88_13_c12 & bh86_w88_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1159_In1_c12 <= "" & bh86_w89_13_c12;
   bh86_w88_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_c12(0);
   bh86_w89_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_c12(1);
   bh86_w90_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1159: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1159_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1159_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_copy1160_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1159_Out0_copy1160_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1161_In0_c12 <= "" & bh86_w90_13_c12 & bh86_w90_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1161_In1_c12 <= "" & bh86_w91_12_c12;
   bh86_w90_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_c12(0);
   bh86_w91_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_c12(1);
   bh86_w92_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1161: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1161_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1161_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_copy1162_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1161_Out0_copy1162_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1163_In0_c12 <= "" & bh86_w92_11_c12 & bh86_w92_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1163_In1_c12 <= "" & bh86_w93_13_c12;
   bh86_w92_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_c12(0);
   bh86_w93_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_c12(1);
   bh86_w94_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1163: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1163_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1163_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_copy1164_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1163_Out0_copy1164_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1165_In0_c12 <= "" & bh86_w95_13_c12 & bh86_w95_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1165_In1_c12 <= "" & bh86_w96_12_c12;
   bh86_w95_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_c12(0);
   bh86_w96_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_c12(1);
   bh86_w97_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1165: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1165_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1165_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_copy1166_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1165_Out0_copy1166_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1167_In0_c12 <= "" & bh86_w97_13_c12 & bh86_w97_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1167_In1_c12 <= "" & bh86_w98_11_c12;
   bh86_w97_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_c12(0);
   bh86_w98_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_c12(1);
   bh86_w99_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1167: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1167_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1167_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_copy1168_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1167_Out0_copy1168_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1169_In0_c12 <= "" & bh86_w99_12_c12 & bh86_w99_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1169_In1_c12 <= "" & bh86_w100_11_c12;
   bh86_w99_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_c12(0);
   bh86_w100_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_c12(1);
   bh86_w101_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1169: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1169_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1169_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_copy1170_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1169_Out0_copy1170_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1171_In0_c12 <= "" & bh86_w101_13_c12 & bh86_w101_14_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1171_In1_c12 <= "" & bh86_w102_10_c12;
   bh86_w101_16_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_c12(0);
   bh86_w102_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_c12(1);
   bh86_w103_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1171: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1171_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1171_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_copy1172_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1171_Out0_copy1172_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1173_In0_c12 <= "" & bh86_w103_12_c12 & bh86_w103_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1173_In1_c12 <= "" & bh86_w104_12_c12;
   bh86_w103_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_c12(0);
   bh86_w104_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_c12(1);
   bh86_w105_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1173: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1173_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1173_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_copy1174_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1173_Out0_copy1174_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1175_In0_c12 <= "" & bh86_w105_11_c12 & bh86_w105_10_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1175_In1_c12 <= "" & bh86_w106_11_c12;
   bh86_w105_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_c12(0);
   bh86_w106_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_c12(1);
   bh86_w107_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1175: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1175_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1175_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_copy1176_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1175_Out0_copy1176_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1177_In0_c12 <= "" & bh86_w107_11_c12 & bh86_w107_10_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1177_In1_c12 <= "" & bh86_w108_11_c12;
   bh86_w107_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_c12(0);
   bh86_w108_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_c12(1);
   bh86_w109_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1177: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1177_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1177_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_copy1178_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1177_Out0_copy1178_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1179_In0_c12 <= "" & bh86_w109_10_c12 & bh86_w109_11_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1179_In1_c12 <= "" & bh86_w110_12_c12;
   bh86_w109_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_c12(0);
   bh86_w110_13_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_c12(1);
   bh86_w111_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1179: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1179_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1179_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_copy1180_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1179_Out0_copy1180_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1181_In0_c12 <= "" & bh86_w112_12_c12 & bh86_w112_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1181_In1_c12 <= "" & bh86_w113_11_c12;
   bh86_w112_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_c12(0);
   bh86_w113_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_c12(1);
   bh86_w114_14_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1181: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1181_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1181_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_copy1182_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1181_Out0_copy1182_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1183_In0_c12 <= "" & bh86_w114_12_c12 & bh86_w114_13_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1183_In1_c12 <= "" & bh86_w115_7_c12;
   bh86_w114_15_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_c12(0);
   bh86_w115_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_c12(1);
   bh86_w116_11_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1183: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1183_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1183_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_copy1184_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1183_Out0_copy1184_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1185_In0_c12 <= "" & bh86_w116_9_c12 & bh86_w116_10_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1185_In1_c12 <= "" & bh86_w117_5_c12;
   bh86_w116_12_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_c12(0);
   bh86_w117_6_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_c12(1);
   bh86_w118_8_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_c12(2);
   Compressor_14_3_Freq300_uid626_uid1185: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1185_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1185_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_copy1186_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1185_Out0_copy1186_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1187_In0_c12 <= "" & bh86_w118_7_c12 & bh86_w118_6_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1187_In1_c12 <= "" & bh86_w119_3_c12;
   bh86_w118_9_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_c12(0);
   bh86_w119_4_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_c12(1);
   Compressor_14_3_Freq300_uid626_uid1187: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1187_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1187_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_copy1188_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_c12 <= Compressor_14_3_Freq300_uid626_bh86_uid1187_Out0_copy1188_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1189_In0_c12 <= "" & bh86_w40_0_c12 & bh86_w40_1_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1189_In1_c12 <= "" & bh86_w41_0_c12 & bh86_w41_1_c12;
   bh86_w40_2_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_c12(0);
   bh86_w41_2_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_c12(1);
   bh86_w42_2_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1189: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1189_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1189_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_copy1190_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1189_Out0_copy1190_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1191_In0_c12 <= "" & bh86_w42_0_c12 & bh86_w42_1_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1191_In1_c12 <= "" & bh86_w43_0_c12 & bh86_w43_1_c12;
   bh86_w42_3_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_c12(0);
   bh86_w43_2_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_c12(1);
   bh86_w44_37_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1191: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1191_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1191_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_copy1192_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1191_Out0_copy1192_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1193_In0_c12 <= "" & bh86_w44_36_c12 & bh86_w44_13_c12 & bh86_w44_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1193_In1_c12 <= "" & bh86_w45_32_c12 & bh86_w45_8_c12;
   bh86_w44_38_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_c12(0);
   bh86_w45_33_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_c12(1);
   bh86_w46_40_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1193: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1193_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1193_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_copy1194_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1193_Out0_copy1194_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1195_In0_c12 <= "" & bh86_w46_39_c12 & bh86_w46_8_c12 & bh86_w46_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1195_In1_c12 <= "" & bh86_w47_43_c12 & bh86_w47_9_c12;
   bh86_w46_41_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_c12(0);
   bh86_w47_44_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_c12(1);
   bh86_w48_46_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_c12(2);
   Compressor_23_3_Freq300_uid650_uid1195: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1195_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1195_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_copy1196_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_c12 <= Compressor_23_3_Freq300_uid650_bh86_uid1195_Out0_copy1196_c12; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1197_In0_c12 <= "" & bh86_w48_45_c12 & bh86_w48_8_c12 & bh86_w48_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1197_In1_c12 <= "" & bh86_w49_46_c12 & bh86_w49_7_c12;
   bh86_w48_47_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_c13(0);
   bh86_w49_47_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_c13(1);
   bh86_w50_46_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1197: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1197_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1197_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_copy1198_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1197_Out0_copy1198_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1199_In0_c12 <= "" & bh86_w50_44_c12 & bh86_w50_45_c12 & bh86_w50_0_c12 & bh86_w50_8_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1199_In1_c12 <= "" & bh86_w51_41_c12;
   bh86_w50_47_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_c13(0);
   bh86_w51_42_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_c13(1);
   bh86_w52_42_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1199: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1199_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1199_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_copy1200_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1199_Out0_copy1200_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1201_In0_c12 <= "" & bh86_w51_0_c12 & bh86_w51_6_c12 & bh86_w51_1_c12;
   bh86_w51_43_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_c12(0);
   bh86_w52_43_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1201: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1201_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_copy1202_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1201_Out0_copy1202_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1203_In0_c12 <= "" & bh86_w52_40_c12 & bh86_w52_41_c12 & bh86_w52_0_c12 & bh86_w52_6_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1203_In1_c12 <= "" & bh86_w53_38_c12;
   bh86_w52_44_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_c13(0);
   bh86_w53_39_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_c13(1);
   bh86_w54_37_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1203: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1203_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1203_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_copy1204_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1203_Out0_copy1204_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1205_In0_c12 <= "" & bh86_w53_0_c12 & bh86_w53_5_c12 & bh86_w53_1_c12;
   bh86_w53_40_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_c12(0);
   bh86_w54_38_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1205: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1205_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_copy1206_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1205_Out0_copy1206_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1207_In0_c12 <= "" & bh86_w54_35_c12 & bh86_w54_36_c12 & bh86_w54_0_c12 & bh86_w54_4_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1207_In1_c12 <= "" & bh86_w55_32_c12;
   bh86_w54_39_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_c13(0);
   bh86_w55_34_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_c13(1);
   bh86_w56_29_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1207: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1207_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1207_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_copy1208_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1207_Out0_copy1208_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1209_In0_c12 <= "" & bh86_w55_33_c12 & bh86_w55_0_c12 & bh86_w55_1_c12 & bh86_w55_3_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1209_In1_c12 <= "" & bh86_w56_28_c12;
   bh86_w55_35_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_c13(0);
   bh86_w56_30_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_c13(1);
   bh86_w57_30_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1209: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1209_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1209_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_copy1210_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1209_Out0_copy1210_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1211_In0_c12 <= "" & bh86_w56_0_c12 & bh86_w56_1_c12 & bh86_w56_3_c12;
   bh86_w56_31_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_c12(0);
   bh86_w57_31_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1211: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1211_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_copy1212_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1211_Out0_copy1212_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1213_In0_c12 <= "" & bh86_w57_28_c12 & bh86_w57_29_c12 & bh86_w57_0_c12 & bh86_w57_1_c12 & bh86_w57_2_c12 & bh86_w57_3_c12;
   bh86_w57_32_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_c13(0);
   bh86_w58_23_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_c13(1);
   bh86_w59_27_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1213: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1213_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_copy1214_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1213_Out0_copy1214_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1215_In0_c12 <= "" & bh86_w58_22_c12 & bh86_w58_0_c12 & bh86_w58_1_c12 & bh86_w58_2_c12 & bh86_w58_3_c12;
   bh86_w58_24_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_c13(0);
   bh86_w59_28_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_c13(1);
   bh86_w60_22_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1215: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1215_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_copy1216_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1215_Out0_copy1216_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1217_In0_c12 <= "" & bh86_w59_25_c12 & bh86_w59_26_c12 & bh86_w59_0_c12 & bh86_w59_1_c12 & bh86_w59_2_c12 & bh86_w59_3_c12;
   bh86_w59_29_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_c13(0);
   bh86_w60_23_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_c13(1);
   bh86_w61_23_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1217: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1217_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_copy1218_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1217_Out0_copy1218_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1219_In0_c12 <= "" & bh86_w60_21_c12 & bh86_w60_0_c12 & bh86_w60_1_c12 & bh86_w60_2_c12 & bh86_w60_3_c12;
   bh86_w60_24_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_c13(0);
   bh86_w61_24_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_c13(1);
   bh86_w62_19_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1219: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1219_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_copy1220_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1219_Out0_copy1220_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1221_In0_c12 <= "" & bh86_w61_21_c12 & bh86_w61_22_c12 & bh86_w61_0_c12 & bh86_w61_1_c12 & bh86_w61_2_c12 & bh86_w61_3_c12;
   bh86_w61_25_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_c13(0);
   bh86_w62_20_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_c13(1);
   bh86_w63_20_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1221: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1221_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_copy1222_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1221_Out0_copy1222_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1223_In0_c12 <= "" & bh86_w62_18_c12 & bh86_w62_0_c12 & bh86_w62_1_c12 & bh86_w62_2_c12 & bh86_w62_3_c12;
   bh86_w62_21_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_c13(0);
   bh86_w63_21_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_c13(1);
   bh86_w64_16_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1223: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1223_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_copy1224_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1223_Out0_copy1224_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1225_In0_c12 <= "" & bh86_w63_18_c12 & bh86_w63_19_c12 & bh86_w63_0_c12 & bh86_w63_1_c12 & bh86_w63_2_c12 & bh86_w63_3_c12;
   bh86_w63_22_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_c13(0);
   bh86_w64_17_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_c13(1);
   bh86_w65_21_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1225: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1225_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_copy1226_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1225_Out0_copy1226_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1227_In0_c12 <= "" & bh86_w64_15_c12 & bh86_w64_0_c12 & bh86_w64_1_c12 & bh86_w64_2_c12 & bh86_w64_3_c12;
   bh86_w64_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_c13(0);
   bh86_w65_22_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_c13(1);
   bh86_w66_14_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1227: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1227_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_copy1228_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1227_Out0_copy1228_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1229_In0_c12 <= "" & bh86_w65_19_c12 & bh86_w65_20_c12 & bh86_w65_0_c12 & bh86_w65_1_c12 & bh86_w65_2_c12 & bh86_w65_3_c12;
   bh86_w65_23_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_c13(0);
   bh86_w66_15_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_c13(1);
   bh86_w67_20_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1229: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1229_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_copy1230_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1229_Out0_copy1230_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1231_In0_c12 <= "" & bh86_w66_13_c12 & bh86_w66_0_c12 & bh86_w66_1_c12 & bh86_w66_2_c12 & bh86_w66_3_c12;
   bh86_w66_16_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_c13(0);
   bh86_w67_21_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_c13(1);
   bh86_w68_15_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1231: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1231_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_copy1232_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1231_Out0_copy1232_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1233_In0_c12 <= "" & bh86_w67_18_c12 & bh86_w67_19_c12 & bh86_w67_0_c12 & bh86_w67_1_c12 & bh86_w67_2_c12 & bh86_w67_3_c12;
   bh86_w67_22_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_c13(0);
   bh86_w68_16_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_c13(1);
   bh86_w69_19_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1233: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1233_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_copy1234_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1233_Out0_copy1234_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1235_In0_c12 <= "" & bh86_w68_14_c12 & bh86_w68_0_c12 & bh86_w68_1_c12 & bh86_w68_2_c12 & bh86_w68_3_c12;
   bh86_w68_17_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_c13(0);
   bh86_w69_20_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_c13(1);
   bh86_w70_17_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1235: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1235_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_copy1236_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1235_Out0_copy1236_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1237_In0_c12 <= "" & bh86_w69_17_c12 & bh86_w69_18_c12 & bh86_w69_0_c12 & bh86_w69_1_c12 & bh86_w69_2_c12 & bh86_w69_3_c12;
   bh86_w69_21_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_c13(0);
   bh86_w70_18_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_c13(1);
   bh86_w71_17_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1237: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1237_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_copy1238_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1237_Out0_copy1238_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1239_In0_c12 <= "" & bh86_w70_16_c12 & bh86_w70_0_c12 & bh86_w70_1_c12 & bh86_w70_2_c12 & bh86_w70_3_c12;
   bh86_w70_19_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_c13(0);
   bh86_w71_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_c13(1);
   bh86_w72_16_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1239: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1239_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_copy1240_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1239_Out0_copy1240_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1241_In0_c12 <= "" & bh86_w71_15_c12 & bh86_w71_0_c12 & bh86_w71_1_c12 & bh86_w71_2_c12 & bh86_w71_3_c12 & bh86_w71_16_c12;
   bh86_w71_19_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_c13(0);
   bh86_w72_17_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_c13(1);
   bh86_w73_17_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1241: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1241_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_copy1242_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1241_Out0_copy1242_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1243_In0_c12 <= "" & bh86_w72_0_c12 & bh86_w72_1_c12 & bh86_w72_2_c12 & bh86_w72_3_c12 & bh86_w72_15_c12;
   bh86_w72_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_c13(0);
   bh86_w73_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_c13(1);
   bh86_w74_16_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1243: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1243_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_copy1244_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1243_Out0_copy1244_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1245_In0_c12 <= "" & bh86_w73_16_c12 & bh86_w73_0_c12 & bh86_w73_1_c12 & bh86_w73_2_c12 & bh86_w73_3_c12 & bh86_w73_15_c12;
   bh86_w73_19_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_c13(0);
   bh86_w74_17_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_c13(1);
   bh86_w75_17_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1245: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1245_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_copy1246_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1245_Out0_copy1246_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1247_In0_c12 <= "" & bh86_w74_15_c12 & bh86_w74_0_c12 & bh86_w74_1_c12 & bh86_w74_2_c12 & bh86_w74_3_c12;
   bh86_w74_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_c13(0);
   bh86_w75_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_c13(1);
   bh86_w76_17_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1247: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1247_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_copy1248_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1247_Out0_copy1248_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1249_In0_c12 <= "" & bh86_w75_15_c12 & bh86_w75_16_c12 & bh86_w75_0_c12 & bh86_w75_1_c12 & bh86_w75_2_c12 & bh86_w75_3_c12;
   bh86_w75_19_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_c13(0);
   bh86_w76_18_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_c13(1);
   bh86_w77_16_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1249: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1249_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_copy1250_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1249_Out0_copy1250_c13; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid958_bh86_uid1251_In0_c12 <= "" & bh86_w76_16_c12 & bh86_w76_0_c12 & bh86_w76_1_c12 & bh86_w76_2_c12 & bh86_w76_3_c12;
   bh86_w76_19_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_c13(0);
   bh86_w77_17_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_c13(1);
   bh86_w78_18_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_c13(2);
   Compressor_5_3_Freq300_uid958_uid1251: Compressor_5_3_Freq300_uid958
      port map ( X0 => Compressor_5_3_Freq300_uid958_bh86_uid1251_In0_c12,
                 R => Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_copy1252_c12);
   Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_c13 <= Compressor_5_3_Freq300_uid958_bh86_uid1251_Out0_copy1252_c13; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1253_In0_c12 <= "" & bh86_w77_14_c12 & bh86_w77_15_c12 & bh86_w77_0_c12 & bh86_w77_1_c12 & bh86_w77_2_c12 & bh86_w77_3_c12;
   bh86_w77_18_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_c13(0);
   bh86_w78_19_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_c13(1);
   bh86_w79_16_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1253: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1253_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_copy1254_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1253_Out0_copy1254_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1255_In0_c12 <= "" & bh86_w78_17_c12 & bh86_w78_0_c12 & bh86_w78_1_c12 & bh86_w78_2_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1255_In1_c12 <= "" & bh86_w79_15_c12;
   bh86_w78_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_c13(0);
   bh86_w79_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_c13(1);
   bh86_w80_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1255: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1255_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1255_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_copy1256_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1255_Out0_copy1256_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1257_In0_c12 <= "" & bh86_w79_0_c12 & bh86_w79_1_c12 & bh86_w79_2_c12;
   bh86_w79_18_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_c12(0);
   bh86_w80_20_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1257: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1257_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_copy1258_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1257_Out0_copy1258_c12; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid616_bh86_uid1259_In0_c12 <= "" & bh86_w80_17_c12 & bh86_w80_18_c12 & bh86_w80_0_c12 & bh86_w80_1_c12 & bh86_w80_2_c12 & bh86_w80_3_c12;
   bh86_w80_21_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_c13(0);
   bh86_w81_15_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_c13(1);
   bh86_w82_18_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_c13(2);
   Compressor_6_3_Freq300_uid616_uid1259: Compressor_6_3_Freq300_uid616
      port map ( X0 => Compressor_6_3_Freq300_uid616_bh86_uid1259_In0_c12,
                 R => Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_copy1260_c12);
   Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_c13 <= Compressor_6_3_Freq300_uid616_bh86_uid1259_Out0_copy1260_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1261_In0_c12 <= "" & bh86_w81_14_c12 & bh86_w81_0_c12 & bh86_w81_1_c12 & bh86_w81_2_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1261_In1_c12 <= "" & bh86_w82_16_c12;
   bh86_w81_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_c13(0);
   bh86_w82_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_c13(1);
   bh86_w83_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1261: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1261_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1261_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_copy1262_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1261_Out0_copy1262_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1263_In0_c12 <= "" & bh86_w82_17_c12 & bh86_w82_0_c12 & bh86_w82_1_c12 & bh86_w82_2_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1263_In1_c12 <= "" & bh86_w83_14_c12;
   bh86_w82_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_c13(0);
   bh86_w83_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_c13(1);
   bh86_w84_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1263: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1263_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1263_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_copy1264_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1263_Out0_copy1264_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1265_In0_c12 <= "" & bh86_w83_0_c12 & bh86_w83_1_c12 & bh86_w83_2_c12;
   bh86_w83_17_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_c12(0);
   bh86_w84_20_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1265: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1265_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_copy1266_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1265_Out0_copy1266_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1267_In0_c12 <= "" & bh86_w84_17_c12 & bh86_w84_18_c12 & bh86_w84_0_c12 & bh86_w84_1_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1267_In1_c12 <= "" & bh86_w85_13_c12;
   bh86_w84_21_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_c13(0);
   bh86_w85_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_c13(1);
   bh86_w86_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1267: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1267_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1267_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_copy1268_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1267_Out0_copy1268_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1269_In0_c12 <= "" & bh86_w85_0_c12 & bh86_w85_1_c12 & bh86_w85_2_c12;
   bh86_w85_15_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_c12(0);
   bh86_w86_19_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1269: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1269_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_copy1270_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1269_Out0_copy1270_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1271_In0_c12 <= "" & bh86_w86_16_c12 & bh86_w86_17_c12 & bh86_w86_0_c12 & bh86_w86_1_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1271_In1_c12 <= "" & bh86_w87_15_c12;
   bh86_w86_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_c13(0);
   bh86_w87_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_c13(1);
   bh86_w88_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1271: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1271_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1271_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_copy1272_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1271_Out0_copy1272_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1273_In0_c12 <= "" & bh86_w87_0_c12 & bh86_w87_1_c12 & bh86_w87_2_c12;
   bh86_w87_17_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_c12(0);
   bh86_w88_17_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_c12(1);
   Compressor_3_2_Freq300_uid712_uid1273: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1273_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_copy1274_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_c12 <= Compressor_3_2_Freq300_uid712_bh86_uid1273_Out0_copy1274_c12; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1275_In0_c12 <= "" & bh86_w88_14_c12 & bh86_w88_0_c12 & bh86_w88_1_c12 & bh86_w88_2_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1275_In1_c12 <= "" & bh86_w89_0_c12;
   bh86_w88_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_c13(0);
   bh86_w89_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_c13(1);
   bh86_w90_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1275: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1275_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1275_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_copy1276_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1275_Out0_copy1276_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1277_In0_c12 <= "" & bh86_w89_1_c12 & bh86_w89_2_c12 & bh86_w89_14_c12;
   bh86_w89_16_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_c13(0);
   bh86_w90_17_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1277: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1277_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_copy1278_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1277_Out0_copy1278_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1279_In0_c12 <= "" & bh86_w90_15_c12 & bh86_w90_0_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1279_In1_c12 <= "" & bh86_w91_13_c12;
   bh86_w90_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_c13(0);
   bh86_w91_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_c13(1);
   bh86_w92_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1279: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1279_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1279_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_copy1280_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1279_Out0_copy1280_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1281_In0_c12 <= "" & bh86_w90_1_c12 & bh86_w90_2_c12 & bh86_w90_14_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1281_In1_c12 <= "" & bh86_w91_0_c12 & bh86_w91_1_c12;
   bh86_w90_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_c13(0);
   bh86_w91_15_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_c13(1);
   bh86_w92_16_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1281: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1281_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1281_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_copy1282_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1281_Out0_copy1282_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1283_In0_c12 <= "" & bh86_w92_13_c12 & bh86_w92_14_c12 & bh86_w92_0_c12 & bh86_w92_1_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c0 <= "" & "0";
   bh86_w92_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_c13(0);
   bh86_w93_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_c13(1);
   bh86_w94_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1283: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1283_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1283_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_copy1284_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1283_Out0_copy1284_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1285_In0_c12 <= "" & bh86_w93_14_c12 & bh86_w93_0_c12 & bh86_w93_1_c12;
   bh86_w93_16_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_c13(0);
   bh86_w94_15_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1285: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1285_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_copy1286_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1285_Out0_copy1286_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1287_In0_c12 <= "" & bh86_w94_12_c12 & bh86_w94_13_c12 & bh86_w94_0_c12 & bh86_w94_1_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c0 <= "" & "0";
   bh86_w94_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_c13(0);
   bh86_w95_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_c13(1);
   bh86_w96_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1287: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1287_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1287_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_copy1288_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1287_Out0_copy1288_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1289_In0_c12 <= "" & bh86_w95_15_c12 & bh86_w95_0_c12 & bh86_w95_1_c12;
   bh86_w95_17_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_c13(0);
   bh86_w96_15_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1289: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1289_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_copy1290_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1289_Out0_copy1290_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1291_In0_c12 <= "" & bh86_w96_13_c12 & bh86_w96_0_c12 & bh86_w96_1_c12;
   bh86_w96_16_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_c13(0);
   bh86_w97_17_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1291: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1291_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_copy1292_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1291_Out0_copy1292_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1293_In0_c12 <= "" & bh86_w97_15_c12 & bh86_w97_16_c12 & bh86_w97_0_c12 & bh86_w97_1_c12;
   Compressor_14_3_Freq300_uid626_bh86_uid1293_In1_c12 <= "" & bh86_w98_12_c12;
   bh86_w97_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_c13(0);
   bh86_w98_13_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_c13(1);
   bh86_w99_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1293: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1293_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1293_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_copy1294_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1293_Out0_copy1294_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1295_In0_c12 <= "" & bh86_w99_14_c12 & bh86_w99_15_c12 & bh86_w99_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1295_In1_c12 <= "" & bh86_w100_12_c12 & bh86_w100_0_c12;
   bh86_w99_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_c13(0);
   bh86_w100_13_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_c13(1);
   bh86_w101_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1295: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1295_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1295_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_copy1296_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1295_Out0_copy1296_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1297_In0_c12 <= "" & bh86_w101_15_c12 & bh86_w101_16_c12 & bh86_w101_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1297_In1_c12 <= "" & bh86_w102_11_c12 & bh86_w102_0_c12;
   bh86_w101_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_c13(0);
   bh86_w102_12_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_c13(1);
   bh86_w103_16_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1297: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1297_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1297_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_copy1298_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1297_Out0_copy1298_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1299_In0_c12 <= "" & bh86_w103_14_c12 & bh86_w103_15_c12 & bh86_w103_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1299_In1_c12 <= "" & bh86_w104_13_c12 & bh86_w104_0_c12;
   bh86_w103_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_c13(0);
   bh86_w104_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_c13(1);
   bh86_w105_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1299: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1299_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1299_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_copy1300_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1299_Out0_copy1300_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1301_In0_c12 <= "" & bh86_w105_12_c12 & bh86_w105_0_c12 & bh86_w105_13_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1301_In1_c12 <= "" & bh86_w106_0_c12 & bh86_w106_12_c12;
   bh86_w105_15_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_c13(0);
   bh86_w106_13_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_c13(1);
   bh86_w107_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1301: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1301_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1301_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_copy1302_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1301_Out0_copy1302_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1303_In0_c12 <= "" & bh86_w107_13_c12 & bh86_w107_0_c12 & bh86_w107_12_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1303_In1_c12 <= "" & bh86_w108_12_c12 & bh86_w108_0_c12;
   bh86_w107_15_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_c13(0);
   bh86_w108_13_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_c13(1);
   bh86_w109_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1303: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1303_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1303_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_copy1304_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1303_Out0_copy1304_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1305_In0_c12 <= "" & bh86_w109_12_c12 & bh86_w109_13_c12 & bh86_w109_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1305_In1_c12 <= "" & bh86_w110_13_c12 & bh86_w110_0_c12;
   bh86_w109_15_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_c13(0);
   bh86_w110_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_c13(1);
   bh86_w111_13_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1305: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1305_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1305_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_copy1306_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1305_Out0_copy1306_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1307_In0_c12 <= "" & bh86_w111_11_c12 & bh86_w111_12_c12 & bh86_w111_0_c12;
   Compressor_23_3_Freq300_uid650_bh86_uid1307_In1_c12 <= "" & bh86_w112_14_c12 & bh86_w112_0_c12;
   bh86_w111_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_c13(0);
   bh86_w112_15_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_c13(1);
   bh86_w113_13_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1307: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1307_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1307_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_copy1308_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1307_Out0_copy1308_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1309_In0_c12 <= "" & bh86_w113_12_c12 & bh86_w113_0_c12 & "0";
   bh86_w113_14_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_c13(0);
   bh86_w114_16_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1309: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1309_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_copy1310_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1309_Out0_copy1310_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1311_In0_c12 <= "" & bh86_w114_14_c12 & bh86_w114_15_c12 & bh86_w114_0_c12;
   bh86_w114_17_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_c13(0);
   bh86_w115_9_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1311: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1311_In0_c12,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_copy1312_c12);
   Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1311_Out0_copy1312_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1313_In0_c12 <= "" & bh86_w116_11_c12 & bh86_w116_12_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1313_In1_c12 <= "" & bh86_w117_6_c12;
   bh86_w116_13_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_c13(0);
   bh86_w117_7_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_c13(1);
   bh86_w118_10_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1313: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1313_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1313_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_copy1314_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1313_Out0_copy1314_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1315_In0_c12 <= "" & bh86_w118_8_c12 & bh86_w118_9_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1315_In1_c12 <= "" & bh86_w119_4_c12;
   bh86_w118_11_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_c13(0);
   bh86_w119_5_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_c13(1);
   Compressor_14_3_Freq300_uid626_uid1315: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1315_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1315_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_copy1316_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1315_Out0_copy1316_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1317_In0_c12 <= "" & bh86_w42_3_c12 & bh86_w42_2_c12 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1317_In1_c12 <= "" & bh86_w43_2_c12;
   bh86_w42_4_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_c13(0);
   bh86_w43_3_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_c13(1);
   bh86_w44_39_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1317: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1317_In0_c12,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1317_In1_c12,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_copy1318_c12);
   Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1317_Out0_copy1318_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1319_In0_c12 <= "" & bh86_w44_38_c12 & bh86_w44_37_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1319_In1_c12 <= "" & bh86_w45_33_c12 & bh86_w45_0_c12;
   bh86_w44_40_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_c13(0);
   bh86_w45_34_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_c13(1);
   bh86_w46_42_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1319: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1319_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1319_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_copy1320_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1319_Out0_copy1320_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1321_In0_c12 <= "" & bh86_w46_40_c12 & bh86_w46_41_c12 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1321_In1_c12 <= "" & bh86_w47_44_c12 & bh86_w47_0_c12;
   bh86_w46_43_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_c13(0);
   bh86_w47_45_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_c13(1);
   bh86_w48_48_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1321: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1321_In0_c12,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1321_In1_c12,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_copy1322_c12);
   Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1321_Out0_copy1322_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1323_In0_c13 <= "" & bh86_w48_46_c13 & bh86_w48_47_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1323_In1_c13 <= "" & bh86_w49_47_c13 & bh86_w49_0_c13;
   bh86_w48_49_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_c13(0);
   bh86_w49_48_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_c13(1);
   bh86_w50_48_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1323: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1323_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1323_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_copy1324_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1323_Out0_copy1324_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1325_In0_c13 <= "" & bh86_w50_46_c13 & bh86_w50_47_c13 & bh86_w50_1_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1325_In1_c13 <= "" & bh86_w51_42_c13 & bh86_w51_43_c13;
   bh86_w50_49_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_c13(0);
   bh86_w51_44_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_c13(1);
   bh86_w52_45_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1325: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1325_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1325_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_copy1326_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1325_Out0_copy1326_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1327_In0_c13 <= "" & bh86_w52_42_c13 & bh86_w52_44_c13 & bh86_w52_1_c13 & bh86_w52_43_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1327_In1_c13 <= "" & bh86_w53_39_c13;
   bh86_w52_46_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_c13(0);
   bh86_w53_41_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_c13(1);
   bh86_w54_40_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1327: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1327_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1327_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_copy1328_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1327_Out0_copy1328_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1329_In0_c13 <= "" & bh86_w54_37_c13 & bh86_w54_39_c13 & bh86_w54_1_c13 & bh86_w54_38_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1329_In1_c13 <= "" & bh86_w55_34_c13;
   bh86_w54_41_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_c13(0);
   bh86_w55_36_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_c13(1);
   bh86_w56_32_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1329: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1329_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1329_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_copy1330_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1329_Out0_copy1330_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1331_In0_c13 <= "" & bh86_w56_29_c13 & bh86_w56_30_c13 & bh86_w56_31_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c0 <= "" & "0" & "0";
   bh86_w56_33_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_c13(0);
   bh86_w57_33_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_c13(1);
   bh86_w58_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1331: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1331_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1331_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_copy1332_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1331_Out0_copy1332_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1333_In0_c13 <= "" & bh86_w57_30_c13 & bh86_w57_32_c13 & bh86_w57_31_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1333_In1_c13 <= "" & bh86_w58_23_c13 & bh86_w58_24_c13;
   bh86_w57_34_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_c13(0);
   bh86_w58_26_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_c13(1);
   bh86_w59_30_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1333: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1333_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1333_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_copy1334_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1333_Out0_copy1334_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1335_In0_c13 <= "" & bh86_w59_27_c13 & bh86_w59_28_c13 & bh86_w59_29_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1335_In1_c13 <= "" & bh86_w60_22_c13 & bh86_w60_23_c13;
   bh86_w59_31_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_c13(0);
   bh86_w60_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_c13(1);
   bh86_w61_26_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1335: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1335_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1335_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_copy1336_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1335_Out0_copy1336_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1337_In0_c13 <= "" & bh86_w61_23_c13 & bh86_w61_24_c13 & bh86_w61_25_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1337_In1_c13 <= "" & bh86_w62_19_c13 & bh86_w62_20_c13;
   bh86_w61_27_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_c13(0);
   bh86_w62_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_c13(1);
   bh86_w63_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1337: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1337_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1337_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_copy1338_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1337_Out0_copy1338_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1339_In0_c13 <= "" & bh86_w63_20_c13 & bh86_w63_21_c13 & bh86_w63_22_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1339_In1_c13 <= "" & bh86_w64_16_c13 & bh86_w64_17_c13;
   bh86_w63_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_c13(0);
   bh86_w64_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_c13(1);
   bh86_w65_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1339: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1339_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1339_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_copy1340_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1339_Out0_copy1340_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1341_In0_c13 <= "" & bh86_w65_21_c13 & bh86_w65_22_c13 & bh86_w65_23_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1341_In1_c13 <= "" & bh86_w66_14_c13 & bh86_w66_15_c13;
   bh86_w65_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_c13(0);
   bh86_w66_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_c13(1);
   bh86_w67_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1341: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1341_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1341_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_copy1342_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1341_Out0_copy1342_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1343_In0_c13 <= "" & bh86_w67_20_c13 & bh86_w67_21_c13 & bh86_w67_22_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1343_In1_c13 <= "" & bh86_w68_15_c13 & bh86_w68_16_c13;
   bh86_w67_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_c13(0);
   bh86_w68_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_c13(1);
   bh86_w69_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1343: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1343_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1343_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_copy1344_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1343_Out0_copy1344_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1345_In0_c13 <= "" & bh86_w69_19_c13 & bh86_w69_20_c13 & bh86_w69_21_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1345_In1_c13 <= "" & bh86_w70_17_c13 & bh86_w70_18_c13;
   bh86_w69_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_c13(0);
   bh86_w70_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_c13(1);
   bh86_w71_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1345: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1345_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1345_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_copy1346_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1345_Out0_copy1346_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1347_In0_c13 <= "" & bh86_w71_17_c13 & bh86_w71_18_c13 & bh86_w71_19_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1347_In1_c13 <= "" & bh86_w72_16_c13 & bh86_w72_17_c13;
   bh86_w71_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_c13(0);
   bh86_w72_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_c13(1);
   bh86_w73_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1347: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1347_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1347_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_copy1348_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1347_Out0_copy1348_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1349_In0_c13 <= "" & bh86_w73_17_c13 & bh86_w73_19_c13 & bh86_w73_18_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1349_In1_c13 <= "" & bh86_w74_17_c13 & bh86_w74_18_c13;
   bh86_w73_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_c13(0);
   bh86_w74_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_c13(1);
   bh86_w75_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1349: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1349_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1349_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_copy1350_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1349_Out0_copy1350_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1351_In0_c13 <= "" & bh86_w75_17_c13 & bh86_w75_18_c13 & bh86_w75_19_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1351_In1_c13 <= "" & bh86_w76_17_c13 & bh86_w76_18_c13;
   bh86_w75_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_c13(0);
   bh86_w76_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_c13(1);
   bh86_w77_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1351: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1351_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1351_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_copy1352_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1351_Out0_copy1352_c13; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid712_bh86_uid1353_In0_c13 <= "" & bh86_w77_16_c13 & bh86_w77_17_c13 & bh86_w77_18_c13;
   bh86_w77_20_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_c13(0);
   bh86_w78_21_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_c13(1);
   Compressor_3_2_Freq300_uid712_uid1353: Compressor_3_2_Freq300_uid712
      port map ( X0 => Compressor_3_2_Freq300_uid712_bh86_uid1353_In0_c13,
                 R => Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_copy1354_c13);
   Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_c13 <= Compressor_3_2_Freq300_uid712_bh86_uid1353_Out0_copy1354_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1355_In0_c13 <= "" & bh86_w78_18_c13 & bh86_w78_19_c13 & bh86_w78_20_c13 & bh86_w78_3_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1355_In1_c13 <= "" & bh86_w79_16_c13;
   bh86_w78_22_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_c13(0);
   bh86_w79_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_c13(1);
   bh86_w80_22_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1355: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1355_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1355_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_copy1356_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1355_Out0_copy1356_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1357_In0_c13 <= "" & bh86_w79_17_c13 & bh86_w79_3_c13 & bh86_w79_18_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c0 <= "" & "0" & "0";
   bh86_w79_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_c13(0);
   bh86_w80_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_c13(1);
   bh86_w81_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1357: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1357_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1357_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_copy1358_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1357_Out0_copy1358_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1359_In0_c13 <= "" & bh86_w80_19_c13 & bh86_w80_21_c13 & bh86_w80_20_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1359_In1_c13 <= "" & bh86_w81_15_c13 & bh86_w81_16_c13;
   bh86_w80_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_c13(0);
   bh86_w81_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_c13(1);
   bh86_w82_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1359: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1359_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1359_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_copy1360_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1359_Out0_copy1360_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1361_In0_c13 <= "" & bh86_w82_18_c13 & bh86_w82_19_c13 & bh86_w82_20_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1361_In1_c13 <= "" & bh86_w83_15_c13 & bh86_w83_16_c13;
   bh86_w82_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_c13(0);
   bh86_w83_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_c13(1);
   bh86_w84_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1361: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1361_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1361_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_copy1362_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1361_Out0_copy1362_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1363_In0_c13 <= "" & bh86_w84_19_c13 & bh86_w84_21_c13 & bh86_w84_2_c13 & bh86_w84_20_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1363_In1_c13 <= "" & bh86_w85_14_c13;
   bh86_w84_23_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_c13(0);
   bh86_w85_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_c13(1);
   bh86_w86_21_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1363: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1363_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1363_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_copy1364_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1363_Out0_copy1364_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1365_In0_c13 <= "" & bh86_w86_18_c13 & bh86_w86_20_c13 & bh86_w86_2_c13 & bh86_w86_19_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1365_In1_c13 <= "" & bh86_w87_16_c13;
   bh86_w86_22_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_c13(0);
   bh86_w87_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_c13(1);
   bh86_w88_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1365: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1365_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1365_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_copy1366_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1365_Out0_copy1366_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1367_In0_c13 <= "" & bh86_w88_16_c13 & bh86_w88_18_c13 & bh86_w88_15_c13 & bh86_w88_17_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1367_In1_c13 <= "" & bh86_w89_15_c13;
   bh86_w88_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_c13(0);
   bh86_w89_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_c13(1);
   bh86_w90_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1367: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1367_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1367_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_copy1368_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1367_Out0_copy1368_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1369_In0_c13 <= "" & bh86_w90_16_c13 & bh86_w90_18_c13 & bh86_w90_19_c13 & bh86_w90_17_c13;
   Compressor_14_3_Freq300_uid626_bh86_uid1369_In1_c13 <= "" & bh86_w91_14_c13;
   bh86_w90_21_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_c13(0);
   bh86_w91_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_c13(1);
   bh86_w92_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1369: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1369_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1369_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_copy1370_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1369_Out0_copy1370_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1371_In0_c13 <= "" & bh86_w92_15_c13 & bh86_w92_17_c13 & bh86_w92_16_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1371_In1_c13 <= "" & bh86_w93_15_c13 & bh86_w93_16_c13;
   bh86_w92_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_c13(0);
   bh86_w93_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_c13(1);
   bh86_w94_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1371: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1371_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1371_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_copy1372_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1371_Out0_copy1372_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1373_In0_c13 <= "" & bh86_w94_14_c13 & bh86_w94_15_c13 & bh86_w94_16_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1373_In1_c13 <= "" & bh86_w95_16_c13 & bh86_w95_17_c13;
   bh86_w94_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_c13(0);
   bh86_w95_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_c13(1);
   bh86_w96_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1373: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1373_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1373_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_copy1374_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1373_Out0_copy1374_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1375_In0_c13 <= "" & bh86_w96_14_c13 & bh86_w96_15_c13 & bh86_w96_16_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1375_In1_c13 <= "" & bh86_w97_17_c13 & bh86_w97_18_c13;
   bh86_w96_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_c13(0);
   bh86_w97_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_c13(1);
   bh86_w98_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1375: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1375_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1375_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_copy1376_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1375_Out0_copy1376_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1377_In0_c13 <= "" & bh86_w98_13_c13 & bh86_w98_0_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1377_In1_c13 <= "" & bh86_w99_16_c13 & bh86_w99_17_c13;
   bh86_w98_15_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_c13(0);
   bh86_w99_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_c13(1);
   bh86_w100_14_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1377: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1377_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1377_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_copy1378_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1377_Out0_copy1378_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1379_In0_c13 <= "" & bh86_w101_17_c13 & bh86_w101_18_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1379_In1_c13 <= "" & bh86_w102_12_c13;
   bh86_w101_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_c13(0);
   bh86_w102_13_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_c13(1);
   bh86_w103_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1379: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1379_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1379_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_copy1380_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1379_Out0_copy1380_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1381_In0_c13 <= "" & bh86_w103_16_c13 & bh86_w103_17_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1381_In1_c13 <= "" & bh86_w104_14_c13;
   bh86_w103_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_c13(0);
   bh86_w104_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_c13(1);
   bh86_w105_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1381: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1381_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1381_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_copy1382_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1381_Out0_copy1382_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1383_In0_c13 <= "" & bh86_w105_14_c13 & bh86_w105_15_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1383_In1_c13 <= "" & bh86_w106_13_c13;
   bh86_w105_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_c13(0);
   bh86_w106_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_c13(1);
   bh86_w107_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1383: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1383_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1383_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_copy1384_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1383_Out0_copy1384_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1385_In0_c13 <= "" & bh86_w107_14_c13 & bh86_w107_15_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1385_In1_c13 <= "" & bh86_w108_13_c13;
   bh86_w107_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_c13(0);
   bh86_w108_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_c13(1);
   bh86_w109_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1385: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1385_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1385_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_copy1386_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1385_Out0_copy1386_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1387_In0_c13 <= "" & bh86_w109_14_c13 & bh86_w109_15_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1387_In1_c13 <= "" & bh86_w110_14_c13;
   bh86_w109_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_c13(0);
   bh86_w110_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_c13(1);
   bh86_w111_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1387: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1387_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1387_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_copy1388_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1387_Out0_copy1388_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1389_In0_c13 <= "" & bh86_w111_13_c13 & bh86_w111_14_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1389_In1_c13 <= "" & bh86_w112_15_c13;
   bh86_w111_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_c13(0);
   bh86_w112_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_c13(1);
   bh86_w113_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1389: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1389_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1389_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_copy1390_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1389_Out0_copy1390_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1391_In0_c13 <= "" & bh86_w113_13_c13 & bh86_w113_14_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1391_In1_c13 <= "" & bh86_w114_16_c13 & bh86_w114_17_c13;
   bh86_w113_16_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_c13(0);
   bh86_w114_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_c13(1);
   bh86_w115_10_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1391: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1391_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1391_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_copy1392_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1391_Out0_copy1392_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1393_In0_c13 <= "" & bh86_w115_8_c13 & bh86_w115_9_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1393_In1_c13 <= "" & bh86_w116_13_c13;
   bh86_w115_11_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_c13(0);
   bh86_w116_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_c13(1);
   bh86_w117_8_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1393: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1393_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1393_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_copy1394_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1393_Out0_copy1394_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1395_In0_c13 <= "" & bh86_w118_10_c13 & bh86_w118_11_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1395_In1_c13 <= "" & bh86_w119_5_c13;
   bh86_w118_12_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_c13(0);
   bh86_w119_6_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_c13(1);
   Compressor_14_3_Freq300_uid626_uid1395: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1395_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1395_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_copy1396_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1395_Out0_copy1396_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1397_In0_c13 <= "" & bh86_w44_40_c13 & bh86_w44_39_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1397_In1_c13 <= "" & bh86_w45_34_c13;
   bh86_w44_41_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_c13(0);
   bh86_w45_35_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_c13(1);
   bh86_w46_44_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1397: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1397_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1397_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_copy1398_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1397_Out0_copy1398_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1399_In0_c13 <= "" & bh86_w46_42_c13 & bh86_w46_43_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1399_In1_c13 <= "" & bh86_w47_45_c13;
   bh86_w46_45_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_c13(0);
   bh86_w47_46_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_c13(1);
   bh86_w48_50_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1399: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1399_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1399_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_copy1400_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1399_Out0_copy1400_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1401_In0_c13 <= "" & bh86_w48_48_c13 & bh86_w48_49_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1401_In1_c13 <= "" & bh86_w49_48_c13;
   bh86_w48_51_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_c13(0);
   bh86_w49_49_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_c13(1);
   bh86_w50_50_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1401: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1401_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1401_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_copy1402_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1401_Out0_copy1402_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1403_In0_c13 <= "" & bh86_w50_48_c13 & bh86_w50_49_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1403_In1_c13 <= "" & bh86_w51_44_c13;
   bh86_w50_51_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_c13(0);
   bh86_w51_45_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_c13(1);
   bh86_w52_47_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1403: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1403_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1403_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_copy1404_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1403_Out0_copy1404_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1405_In0_c13 <= "" & bh86_w52_45_c13 & bh86_w52_46_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1405_In1_c13 <= "" & bh86_w53_41_c13 & bh86_w53_40_c13;
   bh86_w52_48_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_c13(0);
   bh86_w53_42_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_c13(1);
   bh86_w54_42_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1405: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1405_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1405_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_copy1406_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1405_Out0_copy1406_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1407_In0_c13 <= "" & bh86_w54_40_c13 & bh86_w54_41_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1407_In1_c13 <= "" & bh86_w55_35_c13 & bh86_w55_36_c13;
   bh86_w54_43_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_c13(0);
   bh86_w55_37_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_c13(1);
   bh86_w56_34_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1407: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1407_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1407_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_copy1408_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1407_Out0_copy1408_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1409_In0_c13 <= "" & bh86_w56_32_c13 & bh86_w56_33_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1409_In1_c13 <= "" & bh86_w57_33_c13 & bh86_w57_34_c13;
   bh86_w56_35_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_c13(0);
   bh86_w57_35_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_c13(1);
   bh86_w58_27_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1409: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1409_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1409_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_copy1410_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1409_Out0_copy1410_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1411_In0_c13 <= "" & bh86_w58_25_c13 & bh86_w58_26_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1411_In1_c13 <= "" & bh86_w59_30_c13 & bh86_w59_31_c13;
   bh86_w58_28_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_c13(0);
   bh86_w59_32_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_c13(1);
   bh86_w60_26_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1411: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1411_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1411_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_copy1412_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1411_Out0_copy1412_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1413_In0_c13 <= "" & bh86_w60_24_c13 & bh86_w60_25_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1413_In1_c13 <= "" & bh86_w61_26_c13 & bh86_w61_27_c13;
   bh86_w60_27_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_c13(0);
   bh86_w61_28_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_c13(1);
   bh86_w62_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1413: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1413_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1413_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_copy1414_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1413_Out0_copy1414_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1415_In0_c13 <= "" & bh86_w62_21_c13 & bh86_w62_22_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1415_In1_c13 <= "" & bh86_w63_23_c13 & bh86_w63_24_c13;
   bh86_w62_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_c13(0);
   bh86_w63_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_c13(1);
   bh86_w64_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1415: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1415_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1415_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_copy1416_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1415_Out0_copy1416_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1417_In0_c13 <= "" & bh86_w64_18_c13 & bh86_w64_19_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1417_In1_c13 <= "" & bh86_w65_24_c13 & bh86_w65_25_c13;
   bh86_w64_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_c13(0);
   bh86_w65_26_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_c13(1);
   bh86_w66_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1417: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1417_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1417_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_copy1418_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1417_Out0_copy1418_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1419_In0_c13 <= "" & bh86_w66_16_c13 & bh86_w66_17_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1419_In1_c13 <= "" & bh86_w67_23_c13 & bh86_w67_24_c13;
   bh86_w66_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_c13(0);
   bh86_w67_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_c13(1);
   bh86_w68_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1419: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1419_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1419_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_copy1420_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1419_Out0_copy1420_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1421_In0_c13 <= "" & bh86_w68_17_c13 & bh86_w68_18_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1421_In1_c13 <= "" & bh86_w69_22_c13 & bh86_w69_23_c13;
   bh86_w68_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_c13(0);
   bh86_w69_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_c13(1);
   bh86_w70_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1421: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1421_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1421_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_copy1422_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1421_Out0_copy1422_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1423_In0_c13 <= "" & bh86_w70_19_c13 & bh86_w70_20_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1423_In1_c13 <= "" & bh86_w71_20_c13 & bh86_w71_21_c13;
   bh86_w70_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_c13(0);
   bh86_w71_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_c13(1);
   bh86_w72_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1423: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1423_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1423_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_copy1424_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1423_Out0_copy1424_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1425_In0_c13 <= "" & bh86_w72_19_c13 & bh86_w72_18_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1425_In1_c13 <= "" & bh86_w73_20_c13 & bh86_w73_21_c13;
   bh86_w72_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_c13(0);
   bh86_w73_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_c13(1);
   bh86_w74_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1425: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1425_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1425_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_copy1426_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1425_Out0_copy1426_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1427_In0_c13 <= "" & bh86_w74_19_c13 & bh86_w74_16_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1427_In1_c13 <= "" & bh86_w75_20_c13 & bh86_w75_21_c13;
   bh86_w74_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_c13(0);
   bh86_w75_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_c13(1);
   bh86_w76_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1427: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1427_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1427_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_copy1428_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1427_Out0_copy1428_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1429_In0_c13 <= "" & bh86_w76_19_c13 & bh86_w76_20_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1429_In1_c13 <= "" & bh86_w77_19_c13 & bh86_w77_20_c13;
   bh86_w76_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_c13(0);
   bh86_w77_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_c13(1);
   bh86_w78_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1429: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1429_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1429_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_copy1430_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1429_Out0_copy1430_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1431_In0_c13 <= "" & bh86_w78_21_c13 & bh86_w78_22_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1431_In1_c13 <= "" & bh86_w79_19_c13 & bh86_w79_20_c13;
   bh86_w78_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_c13(0);
   bh86_w79_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_c13(1);
   bh86_w80_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1431: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1431_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1431_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_copy1432_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1431_Out0_copy1432_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1433_In0_c13 <= "" & bh86_w80_22_c13 & bh86_w80_23_c13 & bh86_w80_24_c13;
   Compressor_23_3_Freq300_uid650_bh86_uid1433_In1_c13 <= "" & bh86_w81_17_c13 & bh86_w81_18_c13;
   bh86_w80_26_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_c13(0);
   bh86_w81_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_c13(1);
   bh86_w82_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1433: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1433_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1433_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_copy1434_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1433_Out0_copy1434_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1435_In0_c13 <= "" & bh86_w82_21_c13 & bh86_w82_22_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1435_In1_c13 <= "" & bh86_w83_18_c13 & bh86_w83_17_c13;
   bh86_w82_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_c13(0);
   bh86_w83_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_c13(1);
   bh86_w84_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1435: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1435_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1435_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_copy1436_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1435_Out0_copy1436_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1437_In0_c13 <= "" & bh86_w84_22_c13 & bh86_w84_23_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1437_In1_c13 <= "" & bh86_w85_16_c13 & bh86_w85_15_c13;
   bh86_w84_25_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_c13(0);
   bh86_w85_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_c13(1);
   bh86_w86_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1437: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1437_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1437_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_copy1438_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1437_Out0_copy1438_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1439_In0_c13 <= "" & bh86_w86_21_c13 & bh86_w86_22_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1439_In1_c13 <= "" & bh86_w87_18_c13 & bh86_w87_17_c13;
   bh86_w86_24_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_c13(0);
   bh86_w87_19_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_c13(1);
   bh86_w88_21_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1439: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1439_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1439_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_copy1440_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1439_Out0_copy1440_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1441_In0_c13 <= "" & bh86_w88_19_c13 & bh86_w88_20_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1441_In1_c13 <= "" & bh86_w89_17_c13 & bh86_w89_16_c13;
   bh86_w88_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_c13(0);
   bh86_w89_18_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_c13(1);
   bh86_w90_22_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1441: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1441_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1441_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_copy1442_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1441_Out0_copy1442_c13; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid650_bh86_uid1443_In0_c13 <= "" & bh86_w90_20_c13 & bh86_w90_21_c13 & "0";
   Compressor_23_3_Freq300_uid650_bh86_uid1443_In1_c13 <= "" & bh86_w91_16_c13 & bh86_w91_15_c13;
   bh86_w90_23_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_c13(0);
   bh86_w91_17_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_c13(1);
   bh86_w92_20_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_c13(2);
   Compressor_23_3_Freq300_uid650_uid1443: Compressor_23_3_Freq300_uid650
      port map ( X0 => Compressor_23_3_Freq300_uid650_bh86_uid1443_In0_c13,
                 X1 => Compressor_23_3_Freq300_uid650_bh86_uid1443_In1_c13,
                 R => Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_copy1444_c13);
   Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_c13 <= Compressor_23_3_Freq300_uid650_bh86_uid1443_Out0_copy1444_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1445_In0_c13 <= "" & bh86_w92_18_c13 & bh86_w92_19_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1445_In1_c13 <= "" & bh86_w93_17_c13;
   bh86_w92_21_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_c13(0);
   bh86_w93_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_c13(1);
   bh86_w94_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1445: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1445_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1445_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_copy1446_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1445_Out0_copy1446_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1447_In0_c13 <= "" & bh86_w94_17_c13 & bh86_w94_18_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1447_In1_c13 <= "" & bh86_w95_18_c13;
   bh86_w94_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_c13(0);
   bh86_w95_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_c13(1);
   bh86_w96_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1447: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1447_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1447_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_copy1448_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1447_Out0_copy1448_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1449_In0_c13 <= "" & bh86_w96_17_c13 & bh86_w96_18_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1449_In1_c13 <= "" & bh86_w97_19_c13;
   bh86_w96_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_c13(0);
   bh86_w97_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_c13(1);
   bh86_w98_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1449: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1449_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1449_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_copy1450_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1449_Out0_copy1450_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1451_In0_c13 <= "" & bh86_w98_14_c13 & bh86_w98_15_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1451_In1_c13 <= "" & bh86_w99_18_c13;
   bh86_w98_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_c13(0);
   bh86_w99_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_c13(1);
   bh86_w100_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1451: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1451_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1451_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_copy1452_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1451_Out0_copy1452_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1453_In0_c13 <= "" & bh86_w100_13_c13 & bh86_w100_14_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1453_In1_c13 <= "" & bh86_w101_19_c13;
   bh86_w100_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_c13(0);
   bh86_w101_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_c13(1);
   bh86_w102_14_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1453: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1453_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1453_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_copy1454_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1453_Out0_copy1454_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1455_In0_c13 <= "" & bh86_w103_18_c13 & bh86_w103_19_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1455_In1_c13 <= "" & bh86_w104_15_c13;
   bh86_w103_20_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_c13(0);
   bh86_w104_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_c13(1);
   bh86_w105_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1455: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1455_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1455_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_copy1456_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1455_Out0_copy1456_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1457_In0_c13 <= "" & bh86_w105_16_c13 & bh86_w105_17_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1457_In1_c13 <= "" & bh86_w106_14_c13;
   bh86_w105_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_c13(0);
   bh86_w106_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_c13(1);
   bh86_w107_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1457: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1457_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1457_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_copy1458_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1457_Out0_copy1458_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1459_In0_c13 <= "" & bh86_w107_16_c13 & bh86_w107_17_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1459_In1_c13 <= "" & bh86_w108_14_c13;
   bh86_w107_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_c13(0);
   bh86_w108_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_c13(1);
   bh86_w109_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1459: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1459_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1459_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_copy1460_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1459_Out0_copy1460_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1461_In0_c13 <= "" & bh86_w109_16_c13 & bh86_w109_17_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1461_In1_c13 <= "" & bh86_w110_15_c13;
   bh86_w109_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_c13(0);
   bh86_w110_16_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_c13(1);
   bh86_w111_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1461: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1461_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1461_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_copy1462_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1461_Out0_copy1462_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1463_In0_c13 <= "" & bh86_w111_15_c13 & bh86_w111_16_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1463_In1_c13 <= "" & bh86_w112_16_c13;
   bh86_w111_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_c13(0);
   bh86_w112_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_c13(1);
   bh86_w113_17_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1463: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1463_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1463_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_copy1464_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1463_Out0_copy1464_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1465_In0_c13 <= "" & bh86_w113_15_c13 & bh86_w113_16_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1465_In1_c13 <= "" & bh86_w114_18_c13;
   bh86_w113_18_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_c13(0);
   bh86_w114_19_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_c13(1);
   bh86_w115_12_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1465: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1465_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1465_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_copy1466_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1465_Out0_copy1466_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1467_In0_c13 <= "" & bh86_w115_10_c13 & bh86_w115_11_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1467_In1_c13 <= "" & bh86_w116_14_c13;
   bh86_w115_13_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_c13(0);
   bh86_w116_15_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_c13(1);
   bh86_w117_9_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1467: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1467_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1467_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_copy1468_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1467_Out0_copy1468_c13; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid626_bh86_uid1469_In0_c13 <= "" & bh86_w117_7_c13 & bh86_w117_8_c13 & "0" & "0";
   Compressor_14_3_Freq300_uid626_bh86_uid1469_In1_c13 <= "" & bh86_w118_12_c13;
   bh86_w117_10_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_c13(0);
   bh86_w118_13_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_c13(1);
   bh86_w119_7_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_c13(2);
   Compressor_14_3_Freq300_uid626_uid1469: Compressor_14_3_Freq300_uid626
      port map ( X0 => Compressor_14_3_Freq300_uid626_bh86_uid1469_In0_c13,
                 X1 => Compressor_14_3_Freq300_uid626_bh86_uid1469_In1_c13,
                 R => Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_copy1470_c13);
   Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_c13 <= Compressor_14_3_Freq300_uid626_bh86_uid1469_Out0_copy1470_c13; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh86_45_c13 <= bh86_w45_35_c13 & bh86_w44_41_c13 & bh86_w43_3_c13 & bh86_w42_4_c13 & bh86_w41_2_c13 & bh86_w40_2_c13 & bh86_w39_0_c13 & bh86_w38_0_c13 & bh86_w37_0_c13 & bh86_w36_0_c13 & bh86_w35_0_c13 & bh86_w34_0_c13 & bh86_w33_0_c13 & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0";

   bitheapFinalAdd_bh86_In0_c13 <= "0" & bh86_w119_6_c13 & bh86_w118_13_c13 & bh86_w117_9_c13 & bh86_w116_15_c13 & bh86_w115_12_c13 & bh86_w114_19_c13 & bh86_w113_17_c13 & bh86_w112_17_c13 & bh86_w111_17_c13 & bh86_w110_16_c13 & bh86_w109_18_c13 & bh86_w108_15_c13 & bh86_w107_18_c13 & bh86_w106_15_c13 & bh86_w105_18_c13 & bh86_w104_16_c13 & bh86_w103_20_c13 & bh86_w102_13_c13 & bh86_w101_20_c13 & bh86_w100_15_c13 & bh86_w99_19_c13 & bh86_w98_16_c13 & bh86_w97_20_c13 & bh86_w96_19_c13 & bh86_w95_19_c13 & bh86_w94_19_c13 & bh86_w93_18_c13 & bh86_w92_20_c13 & bh86_w91_17_c13 & bh86_w90_22_c13 & bh86_w89_18_c13 & bh86_w88_21_c13 & bh86_w87_19_c13 & bh86_w86_23_c13 & bh86_w85_17_c13 & bh86_w84_24_c13 & bh86_w83_19_c13 & bh86_w82_23_c13 & bh86_w81_19_c13 & bh86_w80_25_c13 & bh86_w79_21_c13 & bh86_w78_23_c13 & bh86_w77_21_c13 & bh86_w76_21_c13 & bh86_w75_22_c13 & bh86_w74_20_c13 & bh86_w73_22_c13 & bh86_w72_20_c13 & bh86_w71_22_c13 & bh86_w70_21_c13 & bh86_w69_24_c13 & bh86_w68_19_c13 & bh86_w67_25_c13 & bh86_w66_18_c13 & bh86_w65_26_c13 & bh86_w64_20_c13 & bh86_w63_25_c13 & bh86_w62_23_c13 & bh86_w61_28_c13 & bh86_w60_26_c13 & bh86_w59_32_c13 & bh86_w58_27_c13 & bh86_w57_35_c13 & bh86_w56_34_c13 & bh86_w55_37_c13 & bh86_w54_42_c13 & bh86_w53_42_c13 & bh86_w52_47_c13 & bh86_w51_45_c13 & bh86_w50_50_c13 & bh86_w49_49_c13 & bh86_w48_50_c13 & bh86_w47_46_c13 & bh86_w46_44_c13;
   bitheapFinalAdd_bh86_In1_c13 <= "0" & bh86_w119_7_c13 & "0" & bh86_w117_10_c13 & "0" & bh86_w115_13_c13 & "0" & bh86_w113_18_c13 & "0" & bh86_w111_18_c13 & "0" & bh86_w109_19_c13 & "0" & bh86_w107_19_c13 & "0" & bh86_w105_19_c13 & "0" & "0" & bh86_w102_14_c13 & "0" & bh86_w100_16_c13 & "0" & bh86_w98_17_c13 & "0" & bh86_w96_20_c13 & "0" & bh86_w94_20_c13 & "0" & bh86_w92_21_c13 & "0" & bh86_w90_23_c13 & "0" & bh86_w88_22_c13 & "0" & bh86_w86_24_c13 & "0" & bh86_w84_25_c13 & "0" & bh86_w82_24_c13 & "0" & bh86_w80_26_c13 & "0" & bh86_w78_24_c13 & "0" & bh86_w76_22_c13 & "0" & bh86_w74_21_c13 & "0" & bh86_w72_21_c13 & "0" & bh86_w70_22_c13 & "0" & bh86_w68_20_c13 & "0" & bh86_w66_19_c13 & "0" & bh86_w64_21_c13 & "0" & bh86_w62_24_c13 & "0" & bh86_w60_27_c13 & "0" & bh86_w58_28_c13 & "0" & bh86_w56_35_c13 & "0" & bh86_w54_43_c13 & "0" & bh86_w52_48_c13 & "0" & bh86_w50_51_c13 & "0" & bh86_w48_51_c13 & "0" & bh86_w46_45_c13;
   bitheapFinalAdd_bh86_Cin_c0 <= '0';

   bitheapFinalAdd_bh86: IntAdder_75_Freq300_uid1472
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 Cin => bitheapFinalAdd_bh86_Cin_c0,
                 X => bitheapFinalAdd_bh86_In0_c13,
                 Y => bitheapFinalAdd_bh86_In1_c13,
                 R => bitheapFinalAdd_bh86_Out_c14);
   bitheapResult_bh86_c14 <= bitheapFinalAdd_bh86_Out_c14(73 downto 0) & tmp_bitheapResult_bh86_45_c14;
   R <= bitheapResult_bh86_c14(119 downto 50);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_80_Freq300_uid1475
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_80_Freq300_uid1475 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
          X : in  std_logic_vector(79 downto 0);
          Y : in  std_logic_vector(79 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(79 downto 0)   );
end entity;

architecture arch of IntAdder_80_Freq300_uid1475 is
signal Rtmp_c14 :  std_logic_vector(79 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11, Y_c12, Y_c13, Y_c14 :  std_logic_vector(79 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Y_c10 <= Y_c9;
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Y_c11 <= Y_c10;
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Y_c12 <= Y_c11;
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Y_c13 <= Y_c12;
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Y_c14 <= Y_c13;
               Cin_c14 <= Cin_c13;
            end if;
         end if;
      end process;
   Rtmp_c14 <= X + Y_c14 + Cin_c14;
   R <= Rtmp_c14;
end architecture;

--------------------------------------------------------------------------------
--                      FPMult_11_66_uid81_Freq300_uid82
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMult_11_66_uid81_Freq300_uid82 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
          X : in  std_logic_vector(11+66+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+67+2 downto 0)   );
end entity;

architecture arch of FPMult_11_66_uid81_Freq300_uid82 is
   component IntMultiplier_67x53_70_Freq300_uid84 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
             X : in  std_logic_vector(66 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(69 downto 0)   );
   end component;

   component IntAdder_80_Freq300_uid1475 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
             X : in  std_logic_vector(79 downto 0);
             Y : in  std_logic_vector(79 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(79 downto 0)   );
   end component;

signal sign_c11, sign_c12, sign_c13, sign_c14 :  std_logic;
signal expX_c11, expX_c12 :  std_logic_vector(10 downto 0);
signal expY_c0, expY_c1, expY_c2, expY_c3, expY_c4, expY_c5, expY_c6, expY_c7, expY_c8, expY_c9, expY_c10, expY_c11, expY_c12 :  std_logic_vector(10 downto 0);
signal expSumPreSub_c12 :  std_logic_vector(12 downto 0);
signal bias_c0, bias_c1, bias_c2, bias_c3, bias_c4, bias_c5, bias_c6, bias_c7, bias_c8, bias_c9, bias_c10, bias_c11, bias_c12 :  std_logic_vector(12 downto 0);
signal expSum_c12, expSum_c13, expSum_c14 :  std_logic_vector(12 downto 0);
signal sigX_c11 :  std_logic_vector(66 downto 0);
signal sigY_c0 :  std_logic_vector(52 downto 0);
signal sigProd_c14 :  std_logic_vector(69 downto 0);
signal excSel_c11 :  std_logic_vector(3 downto 0);
signal exc_c11, exc_c12, exc_c13, exc_c14 :  std_logic_vector(1 downto 0);
signal norm_c14 :  std_logic;
signal expPostNorm_c14 :  std_logic_vector(12 downto 0);
signal sigProdExt_c14 :  std_logic_vector(69 downto 0);
signal expSig_c14 :  std_logic_vector(79 downto 0);
signal round_c0 :  std_logic;
signal expSigPostRound_c14 :  std_logic_vector(79 downto 0);
signal excPostNorm_c14 :  std_logic_vector(1 downto 0);
signal finalExc_c14 :  std_logic_vector(1 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9, Y_c10, Y_c11 :  std_logic_vector(11+52+2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expY_c1 <= expY_c0;
               bias_c1 <= bias_c0;
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               expY_c2 <= expY_c1;
               bias_c2 <= bias_c1;
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               expY_c3 <= expY_c2;
               bias_c3 <= bias_c2;
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               expY_c4 <= expY_c3;
               bias_c4 <= bias_c3;
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               expY_c5 <= expY_c4;
               bias_c5 <= bias_c4;
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               expY_c6 <= expY_c5;
               bias_c6 <= bias_c5;
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               expY_c7 <= expY_c6;
               bias_c7 <= bias_c6;
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               expY_c8 <= expY_c7;
               bias_c8 <= bias_c7;
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               expY_c9 <= expY_c8;
               bias_c9 <= bias_c8;
               Y_c9 <= Y_c8;
            end if;
            if ce_10 = '1' then
               expY_c10 <= expY_c9;
               bias_c10 <= bias_c9;
               Y_c10 <= Y_c9;
            end if;
            if ce_11 = '1' then
               expY_c11 <= expY_c10;
               bias_c11 <= bias_c10;
               Y_c11 <= Y_c10;
            end if;
            if ce_12 = '1' then
               sign_c12 <= sign_c11;
               expX_c12 <= expX_c11;
               expY_c12 <= expY_c11;
               bias_c12 <= bias_c11;
               exc_c12 <= exc_c11;
            end if;
            if ce_13 = '1' then
               sign_c13 <= sign_c12;
               expSum_c13 <= expSum_c12;
               exc_c13 <= exc_c12;
            end if;
            if ce_14 = '1' then
               sign_c14 <= sign_c13;
               expSum_c14 <= expSum_c13;
               exc_c14 <= exc_c13;
            end if;
         end if;
      end process;
   sign_c11 <= X(77) xor Y_c11(63);
   expX_c11 <= X(76 downto 66);
   expY_c0 <= Y(62 downto 52);
   expSumPreSub_c12 <= ("00" & expX_c12) + ("00" & expY_c12);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(1023,13);
   expSum_c12 <= expSumPreSub_c12 - bias_c12;
   sigX_c11 <= "1" & X(65 downto 0);
   sigY_c0 <= "1" & Y(51 downto 0);
   SignificandMultiplication: IntMultiplier_67x53_70_Freq300_uid84
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 X => sigX_c11,
                 Y => sigY_c0,
                 R => sigProd_c14);
   excSel_c11 <= X(79 downto 78) & Y_c11(65 downto 64);
   with excSel_c11  select  
   exc_c11 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c14 <= sigProd_c14(69);
   -- exponent update
   expPostNorm_c14 <= expSum_c14 + ("000000000000" & norm_c14);
   -- significand normalization shift
   sigProdExt_c14 <= sigProd_c14(68 downto 0) & "0" when norm_c14='1' else
                         sigProd_c14(67 downto 0) & "00";
   expSig_c14 <= expPostNorm_c14 & sigProdExt_c14(69 downto 3);
   round_c0 <= '1' ;
   RoundingAdder: IntAdder_80_Freq300_uid1475
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 Cin => round_c0,
                 X => expSig_c14,
                 Y => "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
                 R => expSigPostRound_c14);
   with expSigPostRound_c14(79 downto 78)  select 
   excPostNorm_c14 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c14  select  
   finalExc_c14 <= exc_c14 when  "11"|"10"|"00",
                       excPostNorm_c14 when others; 
   R <= finalExc_c14 & sign_c14 & expSigPostRound_c14(77 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                  LeftShifter68_by_max_65_Freq300_uid1479
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X S
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter68_by_max_65_Freq300_uid1479 is
    port (clk, ce_15, ce_16, ce_17 : in std_logic;
          X : in  std_logic_vector(67 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(132 downto 0)   );
end entity;

architecture arch of LeftShifter68_by_max_65_Freq300_uid1479 is
signal ps_c15, ps_c16, ps_c17 :  std_logic_vector(6 downto 0);
signal level0_c14, level0_c15 :  std_logic_vector(67 downto 0);
signal level1_c15 :  std_logic_vector(68 downto 0);
signal level2_c15 :  std_logic_vector(70 downto 0);
signal level3_c15, level3_c16 :  std_logic_vector(74 downto 0);
signal level4_c16 :  std_logic_vector(82 downto 0);
signal level5_c16, level5_c17 :  std_logic_vector(98 downto 0);
signal level6_c17 :  std_logic_vector(130 downto 0);
signal level7_c17 :  std_logic_vector(194 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_15 = '1' then
               level0_c15 <= level0_c14;
            end if;
            if ce_16 = '1' then
               ps_c16 <= ps_c15;
               level3_c16 <= level3_c15;
            end if;
            if ce_17 = '1' then
               ps_c17 <= ps_c16;
               level5_c17 <= level5_c16;
            end if;
         end if;
      end process;
   ps_c15<= S;
   level0_c14<= X;
   level1_c15<= level0_c15 & (0 downto 0 => '0') when ps_c15(0)= '1' else     (0 downto 0 => '0') & level0_c15;
   level2_c15<= level1_c15 & (1 downto 0 => '0') when ps_c15(1)= '1' else     (1 downto 0 => '0') & level1_c15;
   level3_c15<= level2_c15 & (3 downto 0 => '0') when ps_c15(2)= '1' else     (3 downto 0 => '0') & level2_c15;
   level4_c16<= level3_c16 & (7 downto 0 => '0') when ps_c16(3)= '1' else     (7 downto 0 => '0') & level3_c16;
   level5_c16<= level4_c16 & (15 downto 0 => '0') when ps_c16(4)= '1' else     (15 downto 0 => '0') & level4_c16;
   level6_c17<= level5_c17 & (31 downto 0 => '0') when ps_c17(5)= '1' else     (31 downto 0 => '0') & level5_c17;
   level7_c17<= level6_c17 & (63 downto 0 => '0') when ps_c17(6)= '1' else     (63 downto 0 => '0') & level6_c17;
   R <= level7_c17(132 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_15_Freq300_uid1508
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_15_Freq300_uid1508 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17 : in std_logic;
          X : in  std_logic_vector(14 downto 0);
          Y : in  std_logic_vector(14 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of IntAdder_15_Freq300_uid1508 is
signal Rtmp_c17 :  std_logic_vector(14 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
         end if;
      end process;
   Rtmp_c17 <= X + Y + Cin_c17;
   R <= Rtmp_c17;
end architecture;

--------------------------------------------------------------------------------
--                         FixRealKCM_Freq300_uid1483
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1483 is
    port (clk : in std_logic;
          X : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(10 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1483 is
   component FixRealKCM_Freq300_uid1483_T0_Freq300_uid1486 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(14 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid1483_T1_Freq300_uid1489 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(9 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid1483_T2_Freq300_uid1492 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid1496 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_15_Freq300_uid1508 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17 : in std_logic;
             X : in  std_logic_vector(14 downto 0);
             Y : in  std_logic_vector(14 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(14 downto 0)   );
   end component;

signal FixRealKCM_Freq300_uid1483_A0_c17 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid1483_T0_c17 :  std_logic_vector(14 downto 0);
signal FixRealKCM_Freq300_uid1483_T0_copy1487_c17 :  std_logic_vector(14 downto 0);
signal bh1484_w0_0_c17 :  std_logic;
signal bh1484_w1_0_c17 :  std_logic;
signal bh1484_w2_0_c17 :  std_logic;
signal bh1484_w3_0_c17 :  std_logic;
signal bh1484_w4_0_c17 :  std_logic;
signal bh1484_w5_0_c17 :  std_logic;
signal bh1484_w6_0_c17 :  std_logic;
signal bh1484_w7_0_c17 :  std_logic;
signal bh1484_w8_0_c17 :  std_logic;
signal bh1484_w9_0_c17 :  std_logic;
signal bh1484_w10_0_c17 :  std_logic;
signal bh1484_w11_0_c17 :  std_logic;
signal bh1484_w12_0_c17 :  std_logic;
signal bh1484_w13_0_c17 :  std_logic;
signal bh1484_w14_0_c17 :  std_logic;
signal FixRealKCM_Freq300_uid1483_A1_c17 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid1483_T1_c17 :  std_logic_vector(9 downto 0);
signal FixRealKCM_Freq300_uid1483_T1_copy1490_c17 :  std_logic_vector(9 downto 0);
signal bh1484_w0_1_c17 :  std_logic;
signal bh1484_w1_1_c17 :  std_logic;
signal bh1484_w2_1_c17 :  std_logic;
signal bh1484_w3_1_c17 :  std_logic;
signal bh1484_w4_1_c17 :  std_logic;
signal bh1484_w5_1_c17 :  std_logic;
signal bh1484_w6_1_c17 :  std_logic;
signal bh1484_w7_1_c17 :  std_logic;
signal bh1484_w8_1_c17 :  std_logic;
signal bh1484_w9_1_c17 :  std_logic;
signal FixRealKCM_Freq300_uid1483_A2_c17 :  std_logic_vector(2 downto 0);
signal FixRealKCM_Freq300_uid1483_T2_c17 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid1483_T2_copy1493_c17 :  std_logic_vector(4 downto 0);
signal bh1484_w0_2_c17 :  std_logic;
signal bh1484_w1_2_c17 :  std_logic;
signal bh1484_w2_2_c17 :  std_logic;
signal bh1484_w3_2_c17 :  std_logic;
signal bh1484_w4_2_c17 :  std_logic;
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1497_In0_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1497_In1_c17 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_c17 :  std_logic_vector(2 downto 0);
signal bh1484_w0_3_c17 :  std_logic;
signal bh1484_w1_3_c17 :  std_logic;
signal bh1484_w2_3_c17 :  std_logic;
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_copy1498_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1499_In0_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1499_In1_c17 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_c17 :  std_logic_vector(2 downto 0);
signal bh1484_w2_4_c17 :  std_logic;
signal bh1484_w3_3_c17 :  std_logic;
signal bh1484_w4_3_c17 :  std_logic;
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_copy1500_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1501_In0_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1501_In1_c17 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_c17 :  std_logic_vector(2 downto 0);
signal bh1484_w4_4_c17 :  std_logic;
signal bh1484_w5_2_c17 :  std_logic;
signal bh1484_w6_2_c17 :  std_logic;
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_copy1502_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1503_In0_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1503_In1_c17 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_c17 :  std_logic_vector(2 downto 0);
signal bh1484_w6_3_c17 :  std_logic;
signal bh1484_w7_2_c17 :  std_logic;
signal bh1484_w8_2_c17 :  std_logic;
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_copy1504_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1505_In0_c17 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1505_In1_c17 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_c17 :  std_logic_vector(2 downto 0);
signal bh1484_w8_3_c17 :  std_logic;
signal bh1484_w9_2_c17 :  std_logic;
signal bh1484_w10_1_c17 :  std_logic;
signal Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_copy1506_c17 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh1484_0_c17 :  std_logic_vector(0 downto 0);
signal bitheapFinalAdd_bh1484_In0_c17 :  std_logic_vector(14 downto 0);
signal bitheapFinalAdd_bh1484_In1_c17 :  std_logic_vector(14 downto 0);
signal bitheapFinalAdd_bh1484_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh1484_Out_c17 :  std_logic_vector(14 downto 0);
signal bitheapResult_bh1484_c17 :  std_logic_vector(14 downto 0);
signal OutRes_c17 :  std_logic_vector(14 downto 0);
begin
-- This operator multiplies by 1/log(2)
   FixRealKCM_Freq300_uid1483_A0_c17 <= X(12 downto 8);-- input address  m=9  l=5
   FixRealKCM_Freq300_uid1483_Table0: FixRealKCM_Freq300_uid1483_T0_Freq300_uid1486
      port map ( X => FixRealKCM_Freq300_uid1483_A0_c17,
                 Y => FixRealKCM_Freq300_uid1483_T0_copy1487_c17);
   FixRealKCM_Freq300_uid1483_T0_c17 <= FixRealKCM_Freq300_uid1483_T0_copy1487_c17; -- output copy to hold a pipeline register if needed
   bh1484_w0_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(0);
   bh1484_w1_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(1);
   bh1484_w2_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(2);
   bh1484_w3_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(3);
   bh1484_w4_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(4);
   bh1484_w5_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(5);
   bh1484_w6_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(6);
   bh1484_w7_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(7);
   bh1484_w8_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(8);
   bh1484_w9_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(9);
   bh1484_w10_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(10);
   bh1484_w11_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(11);
   bh1484_w12_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(12);
   bh1484_w13_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(13);
   bh1484_w14_0_c17 <= FixRealKCM_Freq300_uid1483_T0_c17(14);
   FixRealKCM_Freq300_uid1483_A1_c17 <= X(7 downto 3);-- input address  m=4  l=0
   FixRealKCM_Freq300_uid1483_Table1: FixRealKCM_Freq300_uid1483_T1_Freq300_uid1489
      port map ( X => FixRealKCM_Freq300_uid1483_A1_c17,
                 Y => FixRealKCM_Freq300_uid1483_T1_copy1490_c17);
   FixRealKCM_Freq300_uid1483_T1_c17 <= FixRealKCM_Freq300_uid1483_T1_copy1490_c17; -- output copy to hold a pipeline register if needed
   bh1484_w0_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(0);
   bh1484_w1_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(1);
   bh1484_w2_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(2);
   bh1484_w3_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(3);
   bh1484_w4_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(4);
   bh1484_w5_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(5);
   bh1484_w6_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(6);
   bh1484_w7_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(7);
   bh1484_w8_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(8);
   bh1484_w9_1_c17 <= FixRealKCM_Freq300_uid1483_T1_c17(9);
   FixRealKCM_Freq300_uid1483_A2_c17 <= X(2 downto 0);-- input address  m=-1  l=-3
   FixRealKCM_Freq300_uid1483_Table2: FixRealKCM_Freq300_uid1483_T2_Freq300_uid1492
      port map ( X => FixRealKCM_Freq300_uid1483_A2_c17,
                 Y => FixRealKCM_Freq300_uid1483_T2_copy1493_c17);
   FixRealKCM_Freq300_uid1483_T2_c17 <= FixRealKCM_Freq300_uid1483_T2_copy1493_c17; -- output copy to hold a pipeline register if needed
   bh1484_w0_2_c17 <= FixRealKCM_Freq300_uid1483_T2_c17(0);
   bh1484_w1_2_c17 <= FixRealKCM_Freq300_uid1483_T2_c17(1);
   bh1484_w2_2_c17 <= FixRealKCM_Freq300_uid1483_T2_c17(2);
   bh1484_w3_2_c17 <= FixRealKCM_Freq300_uid1483_T2_c17(3);
   bh1484_w4_2_c17 <= FixRealKCM_Freq300_uid1483_T2_c17(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq300_uid1496_bh1484_uid1497_In0_c17 <= "" & bh1484_w0_0_c17 & bh1484_w0_1_c17 & bh1484_w0_2_c17;
   Compressor_23_3_Freq300_uid1496_bh1484_uid1497_In1_c17 <= "" & bh1484_w1_0_c17 & bh1484_w1_1_c17;
   bh1484_w0_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_c17(0);
   bh1484_w1_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_c17(1);
   bh1484_w2_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_c17(2);
   Compressor_23_3_Freq300_uid1496_uid1497: Compressor_23_3_Freq300_uid1496
      port map ( X0 => Compressor_23_3_Freq300_uid1496_bh1484_uid1497_In0_c17,
                 X1 => Compressor_23_3_Freq300_uid1496_bh1484_uid1497_In1_c17,
                 R => Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_copy1498_c17);
   Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1497_Out0_copy1498_c17; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1496_bh1484_uid1499_In0_c17 <= "" & bh1484_w2_0_c17 & bh1484_w2_1_c17 & bh1484_w2_2_c17;
   Compressor_23_3_Freq300_uid1496_bh1484_uid1499_In1_c17 <= "" & bh1484_w3_0_c17 & bh1484_w3_1_c17;
   bh1484_w2_4_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_c17(0);
   bh1484_w3_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_c17(1);
   bh1484_w4_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_c17(2);
   Compressor_23_3_Freq300_uid1496_uid1499: Compressor_23_3_Freq300_uid1496
      port map ( X0 => Compressor_23_3_Freq300_uid1496_bh1484_uid1499_In0_c17,
                 X1 => Compressor_23_3_Freq300_uid1496_bh1484_uid1499_In1_c17,
                 R => Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_copy1500_c17);
   Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1499_Out0_copy1500_c17; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1496_bh1484_uid1501_In0_c17 <= "" & bh1484_w4_0_c17 & bh1484_w4_1_c17 & bh1484_w4_2_c17;
   Compressor_23_3_Freq300_uid1496_bh1484_uid1501_In1_c17 <= "" & bh1484_w5_0_c17 & bh1484_w5_1_c17;
   bh1484_w4_4_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_c17(0);
   bh1484_w5_2_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_c17(1);
   bh1484_w6_2_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_c17(2);
   Compressor_23_3_Freq300_uid1496_uid1501: Compressor_23_3_Freq300_uid1496
      port map ( X0 => Compressor_23_3_Freq300_uid1496_bh1484_uid1501_In0_c17,
                 X1 => Compressor_23_3_Freq300_uid1496_bh1484_uid1501_In1_c17,
                 R => Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_copy1502_c17);
   Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1501_Out0_copy1502_c17; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1496_bh1484_uid1503_In0_c17 <= "" & bh1484_w6_0_c17 & bh1484_w6_1_c17 & "0";
   Compressor_23_3_Freq300_uid1496_bh1484_uid1503_In1_c17 <= "" & bh1484_w7_0_c17 & bh1484_w7_1_c17;
   bh1484_w6_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_c17(0);
   bh1484_w7_2_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_c17(1);
   bh1484_w8_2_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_c17(2);
   Compressor_23_3_Freq300_uid1496_uid1503: Compressor_23_3_Freq300_uid1496
      port map ( X0 => Compressor_23_3_Freq300_uid1496_bh1484_uid1503_In0_c17,
                 X1 => Compressor_23_3_Freq300_uid1496_bh1484_uid1503_In1_c17,
                 R => Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_copy1504_c17);
   Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1503_Out0_copy1504_c17; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1496_bh1484_uid1505_In0_c17 <= "" & bh1484_w8_0_c17 & bh1484_w8_1_c17 & "0";
   Compressor_23_3_Freq300_uid1496_bh1484_uid1505_In1_c17 <= "" & bh1484_w9_0_c17 & bh1484_w9_1_c17;
   bh1484_w8_3_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_c17(0);
   bh1484_w9_2_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_c17(1);
   bh1484_w10_1_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_c17(2);
   Compressor_23_3_Freq300_uid1496_uid1505: Compressor_23_3_Freq300_uid1496
      port map ( X0 => Compressor_23_3_Freq300_uid1496_bh1484_uid1505_In0_c17,
                 X1 => Compressor_23_3_Freq300_uid1496_bh1484_uid1505_In1_c17,
                 R => Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_copy1506_c17);
   Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_c17 <= Compressor_23_3_Freq300_uid1496_bh1484_uid1505_Out0_copy1506_c17; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh1484_0_c17(0) <= bh1484_w0_3_c17;

   bitheapFinalAdd_bh1484_In0_c17 <= "0" & bh1484_w14_0_c17 & bh1484_w13_0_c17 & bh1484_w12_0_c17 & bh1484_w11_0_c17 & bh1484_w10_0_c17 & bh1484_w9_2_c17 & bh1484_w8_2_c17 & bh1484_w7_2_c17 & bh1484_w6_2_c17 & bh1484_w5_2_c17 & bh1484_w4_3_c17 & bh1484_w3_2_c17 & bh1484_w2_3_c17 & bh1484_w1_2_c17;
   bitheapFinalAdd_bh1484_In1_c17 <= "0" & "0" & "0" & "0" & "0" & bh1484_w10_1_c17 & "0" & bh1484_w8_3_c17 & "0" & bh1484_w6_3_c17 & "0" & bh1484_w4_4_c17 & bh1484_w3_3_c17 & bh1484_w2_4_c17 & bh1484_w1_3_c17;
   bitheapFinalAdd_bh1484_Cin_c0 <= '0';

   bitheapFinalAdd_bh1484: IntAdder_15_Freq300_uid1508
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 Cin => bitheapFinalAdd_bh1484_Cin_c0,
                 X => bitheapFinalAdd_bh1484_In0_c17,
                 Y => bitheapFinalAdd_bh1484_In1_c17,
                 R => bitheapFinalAdd_bh1484_Out_c17);
   bitheapResult_bh1484_c17 <= bitheapFinalAdd_bh1484_Out_c17(13 downto 0) & tmp_bitheapResult_bh1484_0_c17;
   OutRes_c17 <= bitheapResult_bh1484_c17(14 downto 0);
   R <= OutRes_c17(14 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_68_Freq300_uid1520
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_68_Freq300_uid1520 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18 : in std_logic;
          X : in  std_logic_vector(67 downto 0);
          Y : in  std_logic_vector(67 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(67 downto 0)   );
end entity;

architecture arch of IntAdder_68_Freq300_uid1520 is
signal Rtmp_c18 :  std_logic_vector(67 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
         end if;
      end process;
   Rtmp_c18 <= X + Y + Cin_c18;
   R <= Rtmp_c18;
end architecture;

--------------------------------------------------------------------------------
--                         FixRealKCM_Freq300_uid1510
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid1510 is
    port (clk, ce_18 : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          R : out  std_logic_vector(66 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid1510 is
   component FixRealKCM_Freq300_uid1510_T0_Freq300_uid1513 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(66 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid1510_T1_Freq300_uid1516 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(61 downto 0)   );
   end component;

   component IntAdder_68_Freq300_uid1520 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18 : in std_logic;
             X : in  std_logic_vector(67 downto 0);
             Y : in  std_logic_vector(67 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(67 downto 0)   );
   end component;

signal FixRealKCM_Freq300_uid1510_A0_c17 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid1510_T0_c18 :  std_logic_vector(66 downto 0);
signal FixRealKCM_Freq300_uid1510_T0_copy1514_c17, FixRealKCM_Freq300_uid1510_T0_copy1514_c18 :  std_logic_vector(66 downto 0);
signal bh1511_w0_0_c18 :  std_logic;
signal bh1511_w1_0_c18 :  std_logic;
signal bh1511_w2_0_c18 :  std_logic;
signal bh1511_w3_0_c18 :  std_logic;
signal bh1511_w4_0_c18 :  std_logic;
signal bh1511_w5_0_c18 :  std_logic;
signal bh1511_w6_0_c18 :  std_logic;
signal bh1511_w7_0_c18 :  std_logic;
signal bh1511_w8_0_c18 :  std_logic;
signal bh1511_w9_0_c18 :  std_logic;
signal bh1511_w10_0_c18 :  std_logic;
signal bh1511_w11_0_c18 :  std_logic;
signal bh1511_w12_0_c18 :  std_logic;
signal bh1511_w13_0_c18 :  std_logic;
signal bh1511_w14_0_c18 :  std_logic;
signal bh1511_w15_0_c18 :  std_logic;
signal bh1511_w16_0_c18 :  std_logic;
signal bh1511_w17_0_c18 :  std_logic;
signal bh1511_w18_0_c18 :  std_logic;
signal bh1511_w19_0_c18 :  std_logic;
signal bh1511_w20_0_c18 :  std_logic;
signal bh1511_w21_0_c18 :  std_logic;
signal bh1511_w22_0_c18 :  std_logic;
signal bh1511_w23_0_c18 :  std_logic;
signal bh1511_w24_0_c18 :  std_logic;
signal bh1511_w25_0_c18 :  std_logic;
signal bh1511_w26_0_c18 :  std_logic;
signal bh1511_w27_0_c18 :  std_logic;
signal bh1511_w28_0_c18 :  std_logic;
signal bh1511_w29_0_c18 :  std_logic;
signal bh1511_w30_0_c18 :  std_logic;
signal bh1511_w31_0_c18 :  std_logic;
signal bh1511_w32_0_c18 :  std_logic;
signal bh1511_w33_0_c18 :  std_logic;
signal bh1511_w34_0_c18 :  std_logic;
signal bh1511_w35_0_c18 :  std_logic;
signal bh1511_w36_0_c18 :  std_logic;
signal bh1511_w37_0_c18 :  std_logic;
signal bh1511_w38_0_c18 :  std_logic;
signal bh1511_w39_0_c18 :  std_logic;
signal bh1511_w40_0_c18 :  std_logic;
signal bh1511_w41_0_c18 :  std_logic;
signal bh1511_w42_0_c18 :  std_logic;
signal bh1511_w43_0_c18 :  std_logic;
signal bh1511_w44_0_c18 :  std_logic;
signal bh1511_w45_0_c18 :  std_logic;
signal bh1511_w46_0_c18 :  std_logic;
signal bh1511_w47_0_c18 :  std_logic;
signal bh1511_w48_0_c18 :  std_logic;
signal bh1511_w49_0_c18 :  std_logic;
signal bh1511_w50_0_c18 :  std_logic;
signal bh1511_w51_0_c18 :  std_logic;
signal bh1511_w52_0_c18 :  std_logic;
signal bh1511_w53_0_c18 :  std_logic;
signal bh1511_w54_0_c18 :  std_logic;
signal bh1511_w55_0_c18 :  std_logic;
signal bh1511_w56_0_c18 :  std_logic;
signal bh1511_w57_0_c18 :  std_logic;
signal bh1511_w58_0_c18 :  std_logic;
signal bh1511_w59_0_c18 :  std_logic;
signal bh1511_w60_0_c18 :  std_logic;
signal bh1511_w61_0_c18 :  std_logic;
signal bh1511_w62_0_c18 :  std_logic;
signal bh1511_w63_0_c18 :  std_logic;
signal bh1511_w64_0_c18 :  std_logic;
signal bh1511_w65_0_c18 :  std_logic;
signal bh1511_w66_0_c18 :  std_logic;
signal FixRealKCM_Freq300_uid1510_A1_c17 :  std_logic_vector(5 downto 0);
signal FixRealKCM_Freq300_uid1510_T1_c18 :  std_logic_vector(61 downto 0);
signal FixRealKCM_Freq300_uid1510_T1_copy1517_c17, FixRealKCM_Freq300_uid1510_T1_copy1517_c18 :  std_logic_vector(61 downto 0);
signal bh1511_w0_1_c18 :  std_logic;
signal bh1511_w1_1_c18 :  std_logic;
signal bh1511_w2_1_c18 :  std_logic;
signal bh1511_w3_1_c18 :  std_logic;
signal bh1511_w4_1_c18 :  std_logic;
signal bh1511_w5_1_c18 :  std_logic;
signal bh1511_w6_1_c18 :  std_logic;
signal bh1511_w7_1_c18 :  std_logic;
signal bh1511_w8_1_c18 :  std_logic;
signal bh1511_w9_1_c18 :  std_logic;
signal bh1511_w10_1_c18 :  std_logic;
signal bh1511_w11_1_c18 :  std_logic;
signal bh1511_w12_1_c18 :  std_logic;
signal bh1511_w13_1_c18 :  std_logic;
signal bh1511_w14_1_c18 :  std_logic;
signal bh1511_w15_1_c18 :  std_logic;
signal bh1511_w16_1_c18 :  std_logic;
signal bh1511_w17_1_c18 :  std_logic;
signal bh1511_w18_1_c18 :  std_logic;
signal bh1511_w19_1_c18 :  std_logic;
signal bh1511_w20_1_c18 :  std_logic;
signal bh1511_w21_1_c18 :  std_logic;
signal bh1511_w22_1_c18 :  std_logic;
signal bh1511_w23_1_c18 :  std_logic;
signal bh1511_w24_1_c18 :  std_logic;
signal bh1511_w25_1_c18 :  std_logic;
signal bh1511_w26_1_c18 :  std_logic;
signal bh1511_w27_1_c18 :  std_logic;
signal bh1511_w28_1_c18 :  std_logic;
signal bh1511_w29_1_c18 :  std_logic;
signal bh1511_w30_1_c18 :  std_logic;
signal bh1511_w31_1_c18 :  std_logic;
signal bh1511_w32_1_c18 :  std_logic;
signal bh1511_w33_1_c18 :  std_logic;
signal bh1511_w34_1_c18 :  std_logic;
signal bh1511_w35_1_c18 :  std_logic;
signal bh1511_w36_1_c18 :  std_logic;
signal bh1511_w37_1_c18 :  std_logic;
signal bh1511_w38_1_c18 :  std_logic;
signal bh1511_w39_1_c18 :  std_logic;
signal bh1511_w40_1_c18 :  std_logic;
signal bh1511_w41_1_c18 :  std_logic;
signal bh1511_w42_1_c18 :  std_logic;
signal bh1511_w43_1_c18 :  std_logic;
signal bh1511_w44_1_c18 :  std_logic;
signal bh1511_w45_1_c18 :  std_logic;
signal bh1511_w46_1_c18 :  std_logic;
signal bh1511_w47_1_c18 :  std_logic;
signal bh1511_w48_1_c18 :  std_logic;
signal bh1511_w49_1_c18 :  std_logic;
signal bh1511_w50_1_c18 :  std_logic;
signal bh1511_w51_1_c18 :  std_logic;
signal bh1511_w52_1_c18 :  std_logic;
signal bh1511_w53_1_c18 :  std_logic;
signal bh1511_w54_1_c18 :  std_logic;
signal bh1511_w55_1_c18 :  std_logic;
signal bh1511_w56_1_c18 :  std_logic;
signal bh1511_w57_1_c18 :  std_logic;
signal bh1511_w58_1_c18 :  std_logic;
signal bh1511_w59_1_c18 :  std_logic;
signal bh1511_w60_1_c18 :  std_logic;
signal bh1511_w61_1_c18 :  std_logic;
signal bitheapFinalAdd_bh1511_In0_c18 :  std_logic_vector(67 downto 0);
signal bitheapFinalAdd_bh1511_In1_c18 :  std_logic_vector(67 downto 0);
signal bitheapFinalAdd_bh1511_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh1511_Out_c18 :  std_logic_vector(67 downto 0);
signal bitheapResult_bh1511_c18 :  std_logic_vector(66 downto 0);
signal OutRes_c18 :  std_logic_vector(66 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_18 = '1' then
               FixRealKCM_Freq300_uid1510_T0_copy1514_c18 <= FixRealKCM_Freq300_uid1510_T0_copy1514_c17;
               FixRealKCM_Freq300_uid1510_T1_copy1517_c18 <= FixRealKCM_Freq300_uid1510_T1_copy1517_c17;
            end if;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq300_uid1510_A0_c17 <= X(10 downto 6);-- input address  m=10  l=6
   FixRealKCM_Freq300_uid1510_Table0: FixRealKCM_Freq300_uid1510_T0_Freq300_uid1513
      port map ( X => FixRealKCM_Freq300_uid1510_A0_c17,
                 Y => FixRealKCM_Freq300_uid1510_T0_copy1514_c17);
   FixRealKCM_Freq300_uid1510_T0_c18 <= FixRealKCM_Freq300_uid1510_T0_copy1514_c18; -- output copy to hold a pipeline register if needed
   bh1511_w0_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(0);
   bh1511_w1_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(1);
   bh1511_w2_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(2);
   bh1511_w3_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(3);
   bh1511_w4_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(4);
   bh1511_w5_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(5);
   bh1511_w6_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(6);
   bh1511_w7_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(7);
   bh1511_w8_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(8);
   bh1511_w9_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(9);
   bh1511_w10_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(10);
   bh1511_w11_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(11);
   bh1511_w12_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(12);
   bh1511_w13_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(13);
   bh1511_w14_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(14);
   bh1511_w15_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(15);
   bh1511_w16_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(16);
   bh1511_w17_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(17);
   bh1511_w18_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(18);
   bh1511_w19_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(19);
   bh1511_w20_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(20);
   bh1511_w21_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(21);
   bh1511_w22_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(22);
   bh1511_w23_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(23);
   bh1511_w24_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(24);
   bh1511_w25_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(25);
   bh1511_w26_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(26);
   bh1511_w27_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(27);
   bh1511_w28_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(28);
   bh1511_w29_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(29);
   bh1511_w30_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(30);
   bh1511_w31_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(31);
   bh1511_w32_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(32);
   bh1511_w33_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(33);
   bh1511_w34_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(34);
   bh1511_w35_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(35);
   bh1511_w36_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(36);
   bh1511_w37_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(37);
   bh1511_w38_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(38);
   bh1511_w39_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(39);
   bh1511_w40_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(40);
   bh1511_w41_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(41);
   bh1511_w42_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(42);
   bh1511_w43_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(43);
   bh1511_w44_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(44);
   bh1511_w45_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(45);
   bh1511_w46_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(46);
   bh1511_w47_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(47);
   bh1511_w48_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(48);
   bh1511_w49_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(49);
   bh1511_w50_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(50);
   bh1511_w51_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(51);
   bh1511_w52_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(52);
   bh1511_w53_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(53);
   bh1511_w54_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(54);
   bh1511_w55_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(55);
   bh1511_w56_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(56);
   bh1511_w57_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(57);
   bh1511_w58_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(58);
   bh1511_w59_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(59);
   bh1511_w60_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(60);
   bh1511_w61_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(61);
   bh1511_w62_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(62);
   bh1511_w63_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(63);
   bh1511_w64_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(64);
   bh1511_w65_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(65);
   bh1511_w66_0_c18 <= FixRealKCM_Freq300_uid1510_T0_c18(66);
   FixRealKCM_Freq300_uid1510_A1_c17 <= X(5 downto 0);-- input address  m=5  l=0
   FixRealKCM_Freq300_uid1510_Table1: FixRealKCM_Freq300_uid1510_T1_Freq300_uid1516
      port map ( X => FixRealKCM_Freq300_uid1510_A1_c17,
                 Y => FixRealKCM_Freq300_uid1510_T1_copy1517_c17);
   FixRealKCM_Freq300_uid1510_T1_c18 <= FixRealKCM_Freq300_uid1510_T1_copy1517_c18; -- output copy to hold a pipeline register if needed
   bh1511_w0_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(0);
   bh1511_w1_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(1);
   bh1511_w2_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(2);
   bh1511_w3_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(3);
   bh1511_w4_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(4);
   bh1511_w5_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(5);
   bh1511_w6_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(6);
   bh1511_w7_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(7);
   bh1511_w8_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(8);
   bh1511_w9_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(9);
   bh1511_w10_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(10);
   bh1511_w11_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(11);
   bh1511_w12_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(12);
   bh1511_w13_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(13);
   bh1511_w14_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(14);
   bh1511_w15_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(15);
   bh1511_w16_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(16);
   bh1511_w17_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(17);
   bh1511_w18_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(18);
   bh1511_w19_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(19);
   bh1511_w20_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(20);
   bh1511_w21_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(21);
   bh1511_w22_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(22);
   bh1511_w23_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(23);
   bh1511_w24_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(24);
   bh1511_w25_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(25);
   bh1511_w26_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(26);
   bh1511_w27_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(27);
   bh1511_w28_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(28);
   bh1511_w29_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(29);
   bh1511_w30_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(30);
   bh1511_w31_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(31);
   bh1511_w32_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(32);
   bh1511_w33_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(33);
   bh1511_w34_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(34);
   bh1511_w35_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(35);
   bh1511_w36_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(36);
   bh1511_w37_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(37);
   bh1511_w38_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(38);
   bh1511_w39_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(39);
   bh1511_w40_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(40);
   bh1511_w41_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(41);
   bh1511_w42_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(42);
   bh1511_w43_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(43);
   bh1511_w44_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(44);
   bh1511_w45_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(45);
   bh1511_w46_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(46);
   bh1511_w47_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(47);
   bh1511_w48_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(48);
   bh1511_w49_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(49);
   bh1511_w50_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(50);
   bh1511_w51_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(51);
   bh1511_w52_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(52);
   bh1511_w53_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(53);
   bh1511_w54_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(54);
   bh1511_w55_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(55);
   bh1511_w56_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(56);
   bh1511_w57_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(57);
   bh1511_w58_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(58);
   bh1511_w59_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(59);
   bh1511_w60_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(60);
   bh1511_w61_1_c18 <= FixRealKCM_Freq300_uid1510_T1_c18(61);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh1511_In0_c18 <= "0" & bh1511_w66_0_c18 & bh1511_w65_0_c18 & bh1511_w64_0_c18 & bh1511_w63_0_c18 & bh1511_w62_0_c18 & bh1511_w61_0_c18 & bh1511_w60_0_c18 & bh1511_w59_0_c18 & bh1511_w58_0_c18 & bh1511_w57_0_c18 & bh1511_w56_0_c18 & bh1511_w55_0_c18 & bh1511_w54_0_c18 & bh1511_w53_0_c18 & bh1511_w52_0_c18 & bh1511_w51_0_c18 & bh1511_w50_0_c18 & bh1511_w49_0_c18 & bh1511_w48_0_c18 & bh1511_w47_0_c18 & bh1511_w46_0_c18 & bh1511_w45_0_c18 & bh1511_w44_0_c18 & bh1511_w43_0_c18 & bh1511_w42_0_c18 & bh1511_w41_0_c18 & bh1511_w40_0_c18 & bh1511_w39_0_c18 & bh1511_w38_0_c18 & bh1511_w37_0_c18 & bh1511_w36_0_c18 & bh1511_w35_0_c18 & bh1511_w34_0_c18 & bh1511_w33_0_c18 & bh1511_w32_0_c18 & bh1511_w31_0_c18 & bh1511_w30_0_c18 & bh1511_w29_0_c18 & bh1511_w28_0_c18 & bh1511_w27_0_c18 & bh1511_w26_0_c18 & bh1511_w25_0_c18 & bh1511_w24_0_c18 & bh1511_w23_0_c18 & bh1511_w22_0_c18 & bh1511_w21_0_c18 & bh1511_w20_0_c18 & bh1511_w19_0_c18 & bh1511_w18_0_c18 & bh1511_w17_0_c18 & bh1511_w16_0_c18 & bh1511_w15_0_c18 & bh1511_w14_0_c18 & bh1511_w13_0_c18 & bh1511_w12_0_c18 & bh1511_w11_0_c18 & bh1511_w10_0_c18 & bh1511_w9_0_c18 & bh1511_w8_0_c18 & bh1511_w7_0_c18 & bh1511_w6_0_c18 & bh1511_w5_0_c18 & bh1511_w4_0_c18 & bh1511_w3_0_c18 & bh1511_w2_0_c18 & bh1511_w1_0_c18 & bh1511_w0_0_c18;
   bitheapFinalAdd_bh1511_In1_c18 <= "0" & "0" & "0" & "0" & "0" & "0" & bh1511_w61_1_c18 & bh1511_w60_1_c18 & bh1511_w59_1_c18 & bh1511_w58_1_c18 & bh1511_w57_1_c18 & bh1511_w56_1_c18 & bh1511_w55_1_c18 & bh1511_w54_1_c18 & bh1511_w53_1_c18 & bh1511_w52_1_c18 & bh1511_w51_1_c18 & bh1511_w50_1_c18 & bh1511_w49_1_c18 & bh1511_w48_1_c18 & bh1511_w47_1_c18 & bh1511_w46_1_c18 & bh1511_w45_1_c18 & bh1511_w44_1_c18 & bh1511_w43_1_c18 & bh1511_w42_1_c18 & bh1511_w41_1_c18 & bh1511_w40_1_c18 & bh1511_w39_1_c18 & bh1511_w38_1_c18 & bh1511_w37_1_c18 & bh1511_w36_1_c18 & bh1511_w35_1_c18 & bh1511_w34_1_c18 & bh1511_w33_1_c18 & bh1511_w32_1_c18 & bh1511_w31_1_c18 & bh1511_w30_1_c18 & bh1511_w29_1_c18 & bh1511_w28_1_c18 & bh1511_w27_1_c18 & bh1511_w26_1_c18 & bh1511_w25_1_c18 & bh1511_w24_1_c18 & bh1511_w23_1_c18 & bh1511_w22_1_c18 & bh1511_w21_1_c18 & bh1511_w20_1_c18 & bh1511_w19_1_c18 & bh1511_w18_1_c18 & bh1511_w17_1_c18 & bh1511_w16_1_c18 & bh1511_w15_1_c18 & bh1511_w14_1_c18 & bh1511_w13_1_c18 & bh1511_w12_1_c18 & bh1511_w11_1_c18 & bh1511_w10_1_c18 & bh1511_w9_1_c18 & bh1511_w8_1_c18 & bh1511_w7_1_c18 & bh1511_w6_1_c18 & bh1511_w5_1_c18 & bh1511_w4_1_c18 & bh1511_w3_1_c18 & bh1511_w2_1_c18 & bh1511_w1_1_c18 & bh1511_w0_1_c18;
   bitheapFinalAdd_bh1511_Cin_c0 <= '0';

   bitheapFinalAdd_bh1511: IntAdder_68_Freq300_uid1520
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 Cin => bitheapFinalAdd_bh1511_Cin_c0,
                 X => bitheapFinalAdd_bh1511_In0_c18,
                 Y => bitheapFinalAdd_bh1511_In1_c18,
                 R => bitheapFinalAdd_bh1511_Out_c18);
   bitheapResult_bh1511_c18 <= bitheapFinalAdd_bh1511_Out_c18(66 downto 0);
   OutRes_c18 <= bitheapResult_bh1511_c18(66 downto 0);
   R <= OutRes_c18(66 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_56_Freq300_uid1523
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_Freq300_uid1523 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19 : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_Freq300_uid1523 is
signal Rtmp_c19 :  std_logic_vector(55 downto 0);
signal X_c18, X_c19 :  std_logic_vector(55 downto 0);
signal Y_c19 :  std_logic_vector(55 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               X_c18 <= X;
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               X_c19 <= X_c18;
               Y_c19 <= Y;
               Cin_c19 <= Cin_c18;
            end if;
         end if;
      end process;
   Rtmp_c19 <= X_c19 + Y_c19 + Cin_c19;
   R <= Rtmp_c19;
end architecture;

--------------------------------------------------------------------------------
--            compressedTable_Freq300_uid1527_diff_Freq300_uid1532
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq300_uid1527_diff_Freq300_uid1532 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of compressedTable_Freq300_uid1527_diff_Freq300_uid1532 is
signal Y0_c19 :  std_logic_vector(49 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c19 :  std_logic_vector(49 downto 0);
begin
   with X  select  Y0_c19 <= 
      "00000000000000000000000000000000000000000000000000" when "0000000000",
      "00010000000000100000000000101010101011010101010110" when "0000000001",
      "00100000000010000000000101010101100000000000010001" when "0000000010",
      "00110000000100100000010010000000110110000010000010" when "0000000011",
      "01000000001000000000101010101101010101011101111000" when "0000000100",
      "01010000001100100001010011011011110110011010000100" when "0000000101",
      "01100000010010000010010000001101100001000000110111" when "0000000110",
      "01110000011000100011100101000011101101100001100011" when "0000000111",
      "00000000100000000101010110000000000100010001011011" when "0000001000",
      "00010000101000100111100111000100011101101100110011" when "0000001001",
      "00100000110010001010011100010011000010011000000010" when "0000001010",
      "00110000111100101101111001101110001011000000100000" when "0000001011",
      "01000001001000010010000011011000100000011101101010" when "0000001100",
      "01010001010100110110111101010100111011110010000000" when "0000001101",
      "01100001100010011100101011100110100110001100000110" when "0000001110",
      "01110001110001000011010010010000111001000111100111" when "0000001111",
      "00000010000000101010110101010111011110001110010001" when "0000010000",
      "00010010010001010011011000111110001111011000111101" when "0000010001",
      "00100010100010111101000001001001010110110000101001" when "0000010010",
      "00110010110101100111110001111101001110101111011110" when "0000010011",
      "01000011001001010011101111011110100010000001101110" when "0000010100",
      "01010011011110000000111101110010001011100110110110" when "0000010101",
      "01100011110011101111100000111101010110110010100001" when "0000010110",
      "01110100001010011111011101000101011111001101101000" when "0000010111",
      "00000100100010010000110110010000010000110111010001" when "0000011000",
      "00010100111011000011110000100011101000000101110110" when "0000011001",
      "00100101010100111000010000000101110001100111111111" when "0000011010",
      "00110101101111101110011000111101001010100101101100" when "0000011011",
      "01000110001011100110001111010000100000100001001111" when "0000011100",
      "01010110101000011111110111000110110001011000010011" when "0000011101",
      "01100111000110011011010100100111001011100100111011" when "0000011110",
      "01110111100101011000101011111001001101111110100101" when "0000011111",
      "00001000000101011000000001000100100111111011001010" when "0000100000",
      "00011000100110011001011000010001011001010000000010" when "0000100001",
      "00101001001000011100110101100111110010010011001000" when "0000100010",
      "00111001101011100010011101010000010011111011110101" when "0000100011",
      "01001010001111101010010011010011101111100100001001" when "0000100100",
      "01011010110100110100011011111011000111001001101011" when "0000100101",
      "01101011011011000000111011001111101101001110101010" when "0000100110",
      "01111100000010001111110101011011000100111011000001" when "0000100111",
      "00001100101010100001001110100111000001111101011000" when "0000101000",
      "00011101010011110101001010111101101000101100001000" when "0000101001",
      "00101101111110001011101110101001001110000110011011" when "0000101010",
      "00111110101001100100111101110100010111110101010011" when "0000101011",
      "01001111010110000000111100101001111100001100100111" when "0000101100",
      "01100000000011011111101111010101000010001100001011" when "0000101101",
      "01110000110010000001011010000001000001100000101111" when "0000101110",
      "10000001100001100110000000111001100010100101000100" when "0000101111",
      "00010010010010001101101000001010011110100010111100" when "0000110000",
      "00100011000011111000010011111111111111010100010011" when "0000110001",
      "00110011110110100110001000100110011111100100001011" when "0000110010",
      "01000100101010010111001010001010101010101111110011" when "0000110011",
      "01010101011111001011011100111001011101000111101001" when "0000110100",
      "01100110010101000011000101000000000011110000100000" when "0000110101",
      "01110111001011111110000110101011111100100100011111" when "0000110110",
      "10001000000011111100100110001010110110010100000101" when "0000110111",
      "00011000111100111110100111101010110000100111010001" when "0000111000",
      "00101001110111000100001111011001111011111110100000" when "0000111001",
      "00111010110010001101100001100110111001110011110100" when "0000111010",
      "01001011101110011010100010100000011100011011110101" when "0000111011",
      "01011100101011101011010110010101100111000110110111" when "0000111100",
      "01101101101010000000000001010101101110000001111101" when "0000111101",
      "01111110101001011000100111110000010110010111111101" when "0000111110",
      "10001111101001110101001101110101010110010010100100" when "0000111111",
      "00100000101011010101110111110100110100111011011000" when "0001000000",
      "00110001101101111010101001111111001010011100111110" when "0001000001",
      "01000010110001100011101000100101000000000100000000" when "0001000010",
      "01010011110110010000110111110111010000000000001100" when "0001000011",
      "01100100111100000010011100000111000101100101011100" when "0001000100",
      "01110110000010111000011001100101111101001100111011" when "0001000101",
      "10000111001010110010110100100101100100010110000100" when "0001000110",
      "10011000010011110001110001010111111001100111101111" when "0001000111",
      "00101001011101110101010100001111001100110001001110" when "0001001000",
      "00111010101000111101100001011101111110101011010011" when "0001001001",
      "01001011110101001010011101010111000001011001011001" when "0001001010",
      "01011101000010011100001100001101011000001010100011" when "0001001011",
      "01101110010000110010110010010100010111011010100101" when "0001001100",
      "01111111100000001110010011111111100100110011000110" when "0001001101",
      "10010000110000101110110101100010110111001100100110" when "0001001110",
      "10100010000010010100011011010010010110101111100101" when "0001001111",
      "00110011010100111111001001100010011100110101100100" when "0001010000",
      "01000100101000101111000100100111110100001010001101" when "0001010001",
      "01010101111101100100010000110111011000101100010110" when "0001010010",
      "01100111010011011110110010100110010111101111001010" when "0001010011",
      "01111000101010011110101110001010001111111011001010" when "0001010100",
      "10001010000010100100000111111000110001001111010101" when "0001010101",
      "10011011011011101111000100000111111101000010001100" when "0001010110",
      "10101100110101111111100111001110000110000010111001" when "0001010111",
      "00111110010001010101110101100001110000011010010011" when "0001011000",
      "01001111101101110001110011011001110001101100000101" when "0001011001",
      "01100001001011010011100101001101010000110111110010" when "0001011010",
      "01110010101001111011001111010011100110011001111110" when "0001011011",
      "10000100001001101000110110000100011100001101010000" when "0001011100",
      "10010101101010011100011101110111101101101011011001" when "0001011101",
      "10100111001100010110001011000101100111101110011101" when "0001011110",
      "10111000101111010110000010000110101000110001110101" when "0001011111",
      "00001010010011011100000111010011100000110011010111" when "0001100000",
      "00011011111000101000011111000101010001010100011011" when "0001100001",
      "00101101011110111011001101110101001101011011000101" when "0001100010",
      "00111111000110010100010111111100111001110011000110" when "0001100011",
      "01010000101110110100000001110110001100101111000110" when "0001100100",
      "01100010011000011010001111111011001110001001101001" when "0001100101",
      "01110100000011000111000110100110010111100110010111" when "0001100110",
      "10000101101110111010101010010010010100010010111111" when "0001100111",
      "00010111011011110100111111011010000001001000100011" when "0001101000",
      "00101001001001110110001010011000101100101100011011" when "0001101001",
      "00111010111000111110001111101001110111010001011100" when "0001101010",
      "01001100101001001101010011101001010010111001000000" when "0001101011",
      "01011110011010100011011010110011000011010100001110" when "0001101100",
      "01110000001101000000101001100011011110000100111101" when "0001101101",
      "10000010000000100101000100010111001010011111000000" when "0001101110",
      "10010011110101010000101111101011000001101001001001" when "0001101111",
      "00100101101011000011101111111100001110011110010100" when "0001110000",
      "00110111100001111110001001101000001101101110101010" when "0001110001",
      "01001001011010000000000001001100101110000000101101" when "0001110010",
      "01011011010011001001011011000111101111110010011011" when "0001110011",
      "01101101001101011010011011110111100101011010011010" when "0001110100",
      "01111111001000110011000111111010110011001000111011" when "0001110101",
      "10010001000101010011100011110000001111001001000110" when "0001110110",
      "10100011000010111011110011110111000001100001111100" when "0001110111",
      "00110101000001101011111100101110100100010111100111" when "0001111000",
      "01000111000001100100000010110110100011101100011010" when "0001111001",
      "01011001000010100100001010101110111101100001111100" when "0001111010",
      "01101011000100101100011000111000000001111010010011" when "0001111011",
      "01111101000111111100110001110010010010111001000110" when "0001111100",
      "10001111001100010101011001111110100100100100101010" when "0001111101",
      "10100001010001110110010101111101111101000111001001" when "0001111110",
      "10110011011000011111101010010001110100101111100111" when "0001111111",
      "00000101100000010001011011011011110101110011010000" when "0010000000",
      "00010111101001001011101101111101111100101110011100" when "0010000001",
      "00101001110011001110100110011010011000000101111011" when "0010000010",
      "00111011111110011010001001010011101000100111111000" when "0010000011",
      "01001110001010101110011011001100100001001101001001" when "0010000100",
      "01100000011000001011100000101000000110111010010011" when "0010000101",
      "01110010100110110001011110001001110001000000110000" when "0010000110",
      "10000100110110100000011000010101001001000000000010" when "0010000111",
      "00010111000111011000010011101110001010100110101111" when "0010001000",
      "00101001011001011001010100111001000011110011110101" when "0010001001",
      "00111011101100100011100000011010010100110111101101" when "0010001010",
      "01001110000000110110111010110110110000010101010100" when "0010001011",
      "01100000010110010011101000110011011011000011011000" when "0010001100",
      "01110010101100111001101110110101101100001101011111" when "0010001101",
      "10000101000100101001010001100011001101010101001110" when "0010001110",
      "10010111011101100010010101100001111010010011011000" when "0010001111",
      "00101001110111100100111111011000000001011001000011" when "0010010000",
      "00111100010010110001010011101100000011010000110001" when "0010010001",
      "01001110101111000111010111000100110010111111101110" when "0010010010",
      "01100001001100100111001110001001010110000110110111" when "0010010011",
      "01110011101011010000111101100001000100100100000011" when "0010010100",
      "10000110001011000100101001110011101000110011001101" when "0010010101",
      "10011000101100000010010111101000111111101111100001" when "0010010110",
      "10101011001110001010001011101001011000110100100011" when "0010010111",
      "00111101110001011100001010011101010101111111010111" when "0010011000",
      "01010000010101111000011000101101101011101111110011" when "0010011001",
      "01100010111011011110111011000011100001001001011111" when "0010011010",
      "01110101100010001111110110001000001111110101000111" when "0010011011",
      "10001000001010001011001110100101100100000001100100" when "0010011100",
      "10011010110011010001001001000101011100100101000010" when "0010011101",
      "10101101011101100001101010010010001010111110001111" when "0010011110",
      "11000000001000111100110110110110010011010101100110" when "0010011111",
      "00010010110101100010110011011100101100011110010101" when "0010100000",
      "00100101100011010011100100110000011111110111101100" when "0010100001",
      "00111000010010001111001111011101001001101110000110" when "0010100010",
      "01001011000010010101111000001110011000111100010101" when "0010100011",
      "01011101110011100111100011110000001111001100101100" when "0010100100",
      "01110000100110000100010110101111000000111010001000" when "0010100101",
      "10000011011001101100010101110111010101010001100000" when "0010100110",
      "10010110001110011111100101110110000110010010101101" when "0010100111",
      "00101001000100011110001011011000100000110001110100" when "0010101000",
      "00111011111011101000001011001100000100011000010100" when "0010101001",
      "01001110110011111101101001111110100011100110010000" when "0010101010",
      "01100001101101011110101100011110000011110011011100" when "0010101011",
      "01110100101000001011010111011000111101010000100101" when "0010101100",
      "10000111100100000011101111011101111011001000100000" when "0010101101",
      "10011010100001000111111001011011111011100001010110" when "0010101110",
      "10101101011111010111111010000010001111011101101011" when "0010101111",
      "00000000011110110011110110000000011010111101110000" when "0010110000",
      "00010011011111011011110010000110010101000000101011" when "0010110001",
      "00100110100001001111110011000100000111100101100011" when "0010110010",
      "00111001100100001111111101101010001111101100101110" when "0010110011",
      "01001100101000011100010110101001011101011000111100" when "0010110100",
      "01011111101101110101000010110010110011110000100100" when "0010110101",
      "01110010110100011010000110110111101000111110101101" when "0010110110",
      "10000101111100001011100111101001100110010100100000" when "0010110111",
      "00011001000101001001101001111010101000001010010000" when "0010111000",
      "00101100001111010100010010011100111110000000100110" when "0010111001",
      "00111111011010101011100110000011001010100001110010" when "0010111010",
      "01010010100111001111101001100000000011100010110101" when "0010111011",
      "01100101110101000000100001100110110010000100101011" when "0010111100",
      "01111001000011111110010011001010110010010101011100" when "0010111101",
      "10001100010100001001000010111111110011110001101001" when "0010111110",
      "10011111100101100000110101111001111001000101010100" when "0010111111",
      "00110010111000000101110000101101011000001101010011" when "0011000000",
      "01000110001011110111111000001110111010011000011001" when "0011000001",
      "01011001100000110111010001010011011100001000100100" when "0011000010",
      "01101100110111000100000000110000001101010100001110" when "0011000011",
      "10000000001110011110001011011010110001000111010010" when "0011000100",
      "10010011100111000101110110001000111110000100100010" when "0011000101",
      "10100111000000111011000101110000111110000110110000" when "0011000110",
      "10111010011011111101111111001001001110100001111101" when "0011000111",
      "00001101111000001110100111001000100000000100100101" when "0011001000",
      "00100001010101101101000010100101110110111000101110" when "0011001001",
      "00110100110100011001010110011000101010100101010111" when "0011001010",
      "01001000010100010011100111011000100110001111100010" when "0011001011",
      "01011011110101011011111010011101101000011011100110" when "0011001100",
      "01101111010111110010010100100000000011001110011011" when "0011001101",
      "10000010111011010110111010011000011100001110100111" when "0011001110",
      "10010110100000001001110000111111101100100101110000" when "0011001111",
      "00101010000110001010111101001111000001000001100110" when "0011010000",
      "00111101101101011010100011111111111001110101010011" when "0011010001",
      "01010001010101111000101010001100001010111010101001" when "0011010010",
      "01100100111111100101010100101101111011110011010100" when "0011010011",
      "01111000101010100000101000011111100111101010000000" when "0011010100",
      "10001100010110101010101010011011111101010011110010" when "0011010101",
      "10100000000100000011011111011101111111010001010000" when "0011010110",
      "10110011110010101011001100100001000011101111101111" when "0011010111",
      "00000111100010100001110110100000110100101010101000" when "0011011000",
      "00011011010011100111100010011001001111101100100001" when "0011011001",
      "00101111000101111100010101000110100110010000011111" when "0011011010",
      "01000010111001100000010011100101011101100011010011" when "0011011011",
      "01010110101110010011100010110010101110100100101101" when "0011011100",
      "01101010100100010110000111101011100110001000100101" when "0011011101",
      "01111110011011101000000111001101100100111000010001" when "0011011110",
      "10010010010100001001100110010110011111010011110000" when "0011011111",
      "00100110001101111010101010000100011101110010111011" when "0011100000",
      "00111010001000111011010111010101111100100110110011" when "0011100001",
      "01001110000101001011110011001001101011111010110101" when "0011100010",
      "01100010000010101100000010011110101111110110000010" when "0011100011",
      "01110110000001011100001010010100100000011100011001" when "0011100100",
      "10001010000001011100001111101010101001101111111011" when "0011100101",
      "10011110000010101100010111100001001011110010000111" when "0011100110",
      "10110010000101001100100110111000011010100100111111" when "0011100111",
      "00000110001000111101000010110000111110001100100001" when "0011101000",
      "00011010001101111101110000001011110010101111110001" when "0011101001",
      "00101110010100001110110100001010001000011010001101" when "0011101010",
      "01000010011011110000010011101101100011011100111011" when "0011101011",
      "01010110100100100010010011110111111100001111111010" when "0011101100",
      "01101010101110100100111001101011011111010011010100" when "0011101101",
      "01111110111001111000001010001010101101010000101101" when "0011101110",
      "10010011000110011100001010011000011010111100010010" when "0011101111",
      "00100111010100010000111111010111110001010110001111" when "0011110000",
      "00111011100011010110101110001100001101101011111001" when "0011110001",
      "01001111110011101101011011111001100001011001000101" when "0011110010",
      "01100100000101010101001101100011110010001001010101" when "0011110011",
      "01111000011000001110001000001111011001111001001010" when "0011110100",
      "10001100101100011000010001000001000110110111010101" when "0011110101",
      "10100001000001110011101100111101111011100110001010" when "0011110110",
      "10110101011000100000100001001011001110111100101111" when "0011110111",
      "00001001110000011110110010101110101100001000001110" when "0011111000",
      "00011110001001101110100110101110010010101101000110" when "0011111001",
      "00110010100100010000000010010000010110101000011111" when "0011111010",
      "01000111000000000011001010011011100000010001010111" when "0011111011",
      "01011011011101001000000100010110101100011001111001" when "0011111100",
      "01101111111011011110110101001001001100010000101001" when "0011111101",
      "10000100011011000111100001111010100101100001111100" when "0011111110",
      "10011000111100000010001111110010110010011001000100" when "0011111111",
      "00101101011110001111000011111010000001100001100110" when "0100000000",
      "01000010000001101110000011011000110110001000101100" when "0100000001",
      "01010110100110011111010011011000000111111110010011" when "0100000010",
      "01101011001100100010111001000001000011010110100010" when "0100000011",
      "01111111110011111000111001011101001001001010111011" when "0100000100",
      "10010100011100100001011001110110001110111011101011" when "0100000101",
      "10101001000110011100011111010110011110110000111111" when "0100000110",
      "10111101110001101010001111001000010111011100010110" when "0100000111",
      "00010010011110001010101110010110101100011001110100" when "0100001000",
      "00100111001011111110000010001100100101110001010100" when "0100001001",
      "00111011111011000100001111110101100000010111111001" when "0100001010",
      "01010000101011011101011100011101001101110001000100" when "0100001011",
      "01100101011101001001101101001111110100010000000111" when "0100001100",
      "01111010010000001001000111011001101110111001010101" when "0100001101",
      "10001111000100011011110000000111101101100011011000" when "0100001110",
      "10100011111010000001101100100110110100111000100010" when "0100001111",
      "00111000110000111011000010000100011110011000000001" when "0100010000",
      "01001101101001000111110101101110011000010111010101" when "0100010001",
      "01100010100010101000001100110010100110000011011101" when "0100010010",
      "01110111011101011100001100011111011111100010010100" when "0100010011",
      "10001100011001100011111010000011110001110011111010" when "0100010100",
      "10100001010110111111011010101110011110110011110000" when "0100010101",
      "10110110010101101110110011101110111101011010000111" when "0100010110",
      "11001011010101110010001010010100111001011101010111" when "0100010111",
      "00100000010111001001100011110000010011110011001111" when "0100011000",
      "00110101011001110101000101010001100010010010001111" when "0100011001",
      "01001010011101110100110100001001001111110010110101" when "0100011010",
      "01011111100011001000110101101000011100010000110110" when "0100011011",
      "01110100101001110001001111000000011100101100110001" when "0100011100",
      "10001001110001101110000101100010111011001101000010" when "0100011101",
      "10011110111010111111011110100001110110111111011011" when "0100011110",
      "10110100000101100101011111001111100100011010010001" when "0100011111",
      "00001001010001100000001100111110101100111101110111" when "0100100000",
      "00011110011110101111101101000010001111010101101111" when "0100100001",
      "00110011101101010100000100101101011111011010000011" when "0100100010",
      "01001000111101001101011001010100000110010000110011" when "0100100011",
      "01011110001110011011110000001010000010001111010000" when "0100100100",
      "01110011100000111111001110100011100110111011001111" when "0100100101",
      "10001000110100110111111001110101011101001100011110" when "0100100110",
      "10011110001010000101110111010100100011001101111000" when "0100100111",
      "00110011100000101001001100010110001100011110111011" when "0100101000",
      "01001000111000100001111110010000000001110101000000" when "0100101001",
      "01011110010001110000010010011000000001011100101100" when "0100101010",
      "01110011101100010100001110000100011110111011001000" when "0100101011",
      "10001001001000001101110110101100000011001111010110" when "0100101100",
      "10011110100101011101010001100101101100110011101000" when "0100101101",
      "10110100000100000010100100001000101111011110110010" when "0100101110",
      "11001001100011111101110011101100110100100101100110" when "0100101111",
      "00011111000101001111000101101001111010111100000010" when "0100110000",
      "00110100100111110110011111011000010110110110101111" when "0100110001",
      "01001010001011110100000110010000110010001100001101" when "0100110010",
      "01011111110001000111111111101100001100010110010011" when "0100110011",
      "01110101010111110010010001000011111010010011011110" when "0100110100",
      "10001010111111110010111111110001100110101000001101" when "0100110101",
      "10100000101001001010010001001111010001100000010001" when "0100110110",
      "10110110010011111000001010110111010000110000001000" when "0100110111",
      "00001011111111111100110010000100001111110110010101" when "0100111000",
      "00100001101101011000001100010001001111111100110010" when "0100111001",
      "00110111011100001010011110111001100111111010001001" when "0100111010",
      "01001101001100010011101111011001000100010011001100" when "0100111011",
      "01100010111101110100000011001011100111011100001001" when "0100111100",
      "01111000110000101011011111101101101001011010000101" when "0100111101",
      "10001110100100111010001010011011111000000100001111" when "0100111110",
      "10100100011010100000001000110011010111000101011010" when "0100111111",
      "00111010010001011101100000010001011111111101010100" when "0101000000",
      "01010000001001110010010110010100000010000001111010" when "0101000001",
      "01100110000011011110110000011001000010100000110110" when "0101000010",
      "01111011111110100010110011111110111100100000110000" when "0101000011",
      "10010001111010111110100110100100100001000010100111" when "0101000100",
      "10100111111000110010001101101000110111000011001110" when "0101000101",
      "10111101110111111101101110101011011011011100011101" when "0101000110",
      "11010011111000100001001111001100000001000110101010" when "0101000111",
      "00101001111010011100110100101010110000111010000111" when "0101001000",
      "00111111111101110000100100101000001001110000010010" when "0101001001",
      "01010110000010011100100100100101000000100101010010" when "0101001010",
      "01101100001000100000111010000010100000011001001100" when "0101001011",
      "10000010001111111101101010100010001010010001100001" when "0101001100",
      "10011000011000110010111011100101110101011010011111" when "0101001101",
      "10101110100011000000110010101111101111001000011111" when "0101001110",
      "11000100101110100111010101100010011010111001011010" when "0101001111",
      "00011010111011100110101001100000110010010110000101" when "0101010000",
      "00110001001001111110110100001110000101010011100110" when "0101010001",
      "01000111011001101111111011001101111001110100110000" when "0101010010",
      "01011101101010111010000100000100001100001011011011" when "0101010011",
      "01110011111101011101010100010101001110111001111100" when "0101010100",
      "10001010010001011001110001100101101010110100011110" when "0101010101",
      "10100000100110101111100001011010011111000010011101" when "0101010110",
      "10110110111101011110101001011001000000111111111101" when "0101010111",
      "00001101010101100111001111000110111100011111000110" when "0101011000",
      "00100011101111001001011000001010010011101001011010" when "0101011001",
      "00111010001010000101001010001001011111000001010010" when "0101011010",
      "01010000100110011010101010101011001101100011010101" when "0101011011",
      "01100111000100001001111111010110100100100111110100" when "0101011100",
      "01111101100011010011001101110011000000000011111111" when "0101011101",
      "10010100000011110110011011101000010010001011100111" when "0101011110",
      "10101010100101110011101110011110100011110010001111" when "0101011111",
      "00000001001001001011001011111110010100001100101101" when "0101100000",
      "00010111101101111100111001110000011001010010100000" when "0101100001",
      "00101110010100001000111101011101111111011111001101" when "0101100010",
      "01000100111011101111011100110000101001110011110110" when "0101100011",
      "01011011100100110000011101010010010001111000011000" when "0101100100",
      "01110010001111001100000100101101000111111101000001" when "0101100101",
      "10001000111011000010011000101011110010111011110010" when "0101100110",
      "10011111101000010011011110111001010000011001110001" when "0101100111",
      "00110110010110111111011101000000110100101000101000" when "0101101000",
      "01001101000111000110011000101110001010101000000010" when "0101101001",
      "01100011111000101000010111101101010100000111000001" when "0101101010",
      "01111010101011100101011111101010101001100101011100" when "0101101011",
      "10010001011111111101110110010010111010010101011011" when "0101101100",
      "10101000010101110001100001010011001100011100110000" when "0101101101",
      "10111111001101000000100110011000111100110110010001" when "0101101110",
      "11010110000101101011001011010001111111010011011000" when "0101101111",
      "00101100111111110001010101101100011110011101011011" when "0101110000",
      "01000011111011010011001011010110111011110111001001" when "0101110001",
      "01011010111000010000110010000000001111111110000010" when "0101110010",
      "01110001110110101010001111010111101010001011111010" when "0101110011",
      "10001000110110011111101001001100110000111000001110" when "0101110100",
      "10011111110111110001000101001111100001011001100010" when "0101110101",
      "10110110111010011110101001010000010000000111000000" when "0101110110",
      "11001101111110101000011010111111101000011001101111" when "0101110111",
      "00100101000100001110100000001110101100101110010011" when "0101111000",
      "00111100001011010000111110101110110110100110000110" when "0101111001",
      "01010011010011101111111100010001110110101000111001" when "0101111010",
      "01101010011101101011011110101001110100100110001101" when "0101111011",
      "10000001101001000011101011101001001111010110101110" when "0101111100",
      "10011000110101111000101001000010111100111101110101" when "0101111101",
      "10110000000100001010011100101010001010101010111111" when "0101111110",
      "11000111010011111001001100010010011100111011001111" when "0101111111",
      "00011110100101000100111101101111101111011010100110" when "0110000000",
      "00110101110111101101110110110110010101000101100011" when "0110000001",
      "01001101001011110011111101011010111000001010100000" when "0110000010",
      "01100100100001010111010111010010011010001011001101" when "0110000011",
      "01111011111000011000001010010010010011111110010000" when "0110000100",
      "10010011010000110110011100010000010101110000100001" when "0110000101",
      "10101010101010110010010011000010100111000110100111" when "0110000110",
      "11000010000110001011110100011111100110111110010111" when "0110000111",
      "00011001100011000011000110011110001011110000001111" when "0110001000",
      "00110001000001011000001110110101100011010000110111" when "0110001001",
      "01001000100001001011010011011101010010110010011101" when "0110001010",
      "01100000000010011100011010001101010111000110010011" when "0110001011",
      "01110111100101001011101000111110000100011110001100" when "0110001100",
      "10001111001001011001000101101000000110101101111100" when "0110001101",
      "10100110101111000100110110000100100001001100110110" when "0110001110",
      "10111110010110001111000000001100101110110111001001" when "0110001111",
      "00010101111110110111101001111010100010001111011110" when "0110010000",
      "00101101101000111110111001001000000101100000011010" when "0110010001",
      "01000101010100100100110011101111111010011101110110" when "0110010010",
      "01011101000001101001011111101100111010100110100110" when "0110010011",
      "01110100110000001101000010111010010111000101110000" when "0110010100",
      "10001100100000001111100011010011111000110100001111" when "0110010101",
      "10100100010001110001000110110101100000011010010010" when "0110010110",
      "10111100000100110001110011011011100110010000111010" when "0110010111",
      "00010011111001010001101111000010111010100011010111" when "0110011000",
      "00101011101111010000111111101000100101010000101011" when "0110011001",
      "01000011100110101111101011001010000110001101001000" when "0110011010",
      "01011011011111101101110111100101010101000011101110" when "0110011011",
      "01110011011010001011101010111000100001010111101100" when "0110011100",
      "10001011010110001001001011000010010010100101111111" when "0110011101",
      "10100011010011100110011110000001101000000110110000" when "0110011110",
      "10111011010010100011101001110101111001001110111000" when "0110011111",
      "00010011010011000000110100011110110101010001011101" when "0110100000",
      "00101011010100111110000011111100100011100001001111" when "0110100001",
      "01000011011000011011011110001111100011010010001111" when "0110100010",
      "01011011011101011001001001011000101011111011001010" when "0110100011",
      "01110011100011110111001011011001001100110110111001" when "0110100100",
      "10001011101011110101101010010010101101100110000100" when "0110100101",
      "10100011110101010100101100000111001101110000100011" when "0110100110",
      "10111100000000010100010110111001000101000110111011" when "0110100111",
      "00010100001100110100110000101011000011100011111111" when "0110101000",
      "00101100011010110101111111100000010001001110010101" when "0110101001",
      "01000100101010011000001001011100001110011001110010" when "0110101010",
      "01011100111011011011010100100010110011101000111101" when "0110101011",
      "01110101001101111111100110111000010001101110101111" when "0110101100",
      "10001101100010000101000110100001010001101111110111" when "0110101101",
      "10100101110111101011111001100010110101000100010110" when "0110101110",
      "10111110001110110100000110000010010101011001000101" when "0110101111",
      "00010110100111011101110010000101100100110001010100" when "0110110000",
      "00101111000001101001000011110010101101101000001100" when "0110110001",
      "01000111011101010110000001010000010010110010010000" when "0110110010",
      "01011111111010100100110000100101001111011111000001" when "0110110011",
      "01111000011001010101010111111000110111011010011010" when "0110110100",
      "10010000111001100111111101010010110110101110011010" when "0110110101",
      "10101001011011011100100110111011010010000100011111" when "0110110110",
      "11000001111110110011011010111010100110100111001011" when "0110110111",
      "00011010100011101100011111011001101010000011100111" when "0110111000",
      "00110011001010000111111010100001101010101011000001" when "0110111001",
      "01001011110010000101110010011100001111010100010110" when "0110111010",
      "01100100011011100110001101010011010111011101101010" when "0110111011",
      "01111101000110101001010001010001011011001101110101" when "0110111100",
      "10010101110011001111000100100001001011010101111110" when "0110111101",
      "10101110100001010111101101001101110001010011000001" when "0110111110",
      "11000111010001000011010001100010101111001111010010" when "0110111111",
      "00100000000010010001110111101100000000000011111110" when "0111000000",
      "00111000110101000011100101110101110111011010101111" when "0111000001",
      "01010001101001011000100010001101000001101111010001" when "0111000010",
      "01101010011111010000110010111110100100010000110010" when "0111000011",
      "10000011010110101100011110010111111101000011100101" when "0111000100",
      "10011100001111101011101010100111000011000010101011" when "0111000101",
      "10110101001010001110011101111010000110000001001110" when "0111000110",
      "11001110000110010100111110011111101110101100001100" when "0111000111",
      "00100111000011111111010010100110111110101011110111" when "0111001000",
      "01000000000011001101100000011111010000100101011000" when "0111001001",
      "01011001000011111111101110011000010111111100010111" when "0111001010",
      "01110010000110010110000010100010100001010100011001" when "0111001011",
      "10001011001010010000100011001110010010010010101010" when "0111001100",
      "10100100001111101111010110101100101001011111011110" when "0111001101",
      "10111101010110110010100011001110111110100111110010" when "0111001110",
      "11010110011111011010001111000111000010011110111010" when "0111001111",
      "00101111101001100110100000100110111110111111111011" when "0111010000",
      "01001000110101010111011110000001010111001111010110" when "0111010001",
      "01100010000010101101001101101001000111011100101010" when "0111010010",
      "01111011010001100111110101110001100101000011111000" when "0111010011",
      "10010100100010000111011100101110011110101111001100" when "0111010100",
      "10101101110100001100001000110011111100011000011101" when "0111010101",
      "11000111000111110110000000010110011111001010110100" when "0111010110",
      "11100000011101000101001001101011000001100100010100" when "0111010111",
      "00111001110011111001101011000110110111010111011010" when "0111011000",
      "01010011001100010011101010111111101101101100100100" when "0111011001",
      "01101100100110010011001111101011101011000011111010" when "0111011010",
      "10000110000001111000011111100001001111010110101111" when "0111011011",
      "10011111011111000011100000110111010011111001001010" when "0111011100",
      "10111000111101110100011010000101001011011011100111" when "0111011101",
      "11010010011110001011010001100010100010001100100011" when "0111011110",
      "11101100000000001000001101100111011101111001111110" when "0111011111",
      "00000101100011101011010100101100011101110011000001" when "0111100000",
      "00011111001000110100101101001010011010101001100111" when "0111100001",
      "00111000101111100100011101011010100110110011111111" when "0111100010",
      "01010010010111111010101011110110101110001110010110" when "0111100011",
      "01101100000001110111011110111000110110011100011011" when "0111100100",
      "10000101101101011010111100111011011110101011001000" when "0111100101",
      "10011111011010100101001100011001011111110010000110" when "0111100110",
      "10111001001001010110010011101110001100010101010101" when "0111100111",
      "00010010111001101110011001010101010000100110110010" when "0111101000",
      "00101100101011101101100011101010110010101000000000" when "0111101001",
      "01000110011111010011111001001011010010001011101101" when "0111101010",
      "01100000010100100001100000010011101000110111011010" when "0111101011",
      "01111010001011010110011111100001001010000101000001" when "0111101100",
      "10010100000011110010111101010001100011000100011110" when "0111101101",
      "10101101111101110111000000000010111010111101010111" when "0111101110",
      "11000111111001100010101110010011110010110000100000" when "0111101111",
      "00100001110110110110001110100011000101011001100101" when "0111110000",
      "00111011110101110001100111010000000111110000110100" when "0111110001",
      "01010101110110010100111110111010101000101100100000" when "0111110010",
      "01101111111000100000011100000010110001000010101101" when "0111110011",
      "10001001111100010100000101001001000011101010110101" when "0111110100",
      "10100100000001110000000000101110011101011111010011" when "0111110101",
      "10111110001000110100010101010100010101011111001000" when "0111110110",
      "11011000010001100001001001011100011100101111100111" when "0111110111",
      "00110010011011110110100011101000111110011101111011" when "0111111000",
      "01001100100111110100101010011100100000000000101111" when "0111111001",
      "01100110110101011011100100011010000000111001111001" when "0111111010",
      "10000001000100101011011000000100111010111000000001" when "0111111011",
      "10011011010101100100001100000001000001111000001011" when "0111111100",
      "10110101101000000110000110110010100100000111011110" when "0111111101",
      "11001111111100010001001110111110001010000100101111" when "0111111110",
      "11101010010010000101101011001000110110100010001011" when "0111111111",
      "00010001011001011111100011011111001011000001010000" when "1000000000",
      "00011011000110111000100100000010011101100011001011" when "1000000001",
      "00100100110100111000011011010111011111000001111011" when "1000000010",
      "00101110100011011111001011111001101111011011010111" when "1000000011",
      "00111000010010101100111000000100111000011011101100" when "1000000100",
      "01000010000010100001100010010100101101011101111111" when "1000000101",
      "01001011110010111101001101000101001011101100111001" when "1000000110",
      "01010101100011111111111010110010011010000011000111" when "1000000111",
      "00011111010101101001101101111000101001001100001010" when "1000001000",
      "00101001000111111010101000110100010011100100110101" when "1000001001",
      "00110010111010110010101110000001111101011011111010" when "1000001010",
      "00111100101110010001111111111110010100110010110010" when "1000001011",
      "01000110100010011000100001000110010001011101111101" when "1000001100",
      "01010000010111000110010011110110110101000101110001" when "1000001101",
      "01011010001100011011011010101101001011000110111110" when "1000001110",
      "01100100000010010111111000000110101000110011010100" when "1000001111",
      "00101101111000111011101110100000101101010010001101" when "1000010000",
      "00110111110000000111000000011001000001100001010010" when "1000010001",
      "01000001100111111001110000001101011000010101000110" when "1000010010",
      "01001011100000010100000000011011101110011001101001" when "1000010011",
      "01010101011001010101110011100010001010010011000001" when "1000010100",
      "01011111010010111111001011111110111100011110000011" when "1000010101",
      "01101001001101010000001100010000011111010000111010" when "1000010110",
      "01110011001000001000110110110101010110111011101110" when "1000010111",
      "00111101000011101001001110001100010001101001001011" when "1000011000",
      "01000110111111110001010100110100000111011111001010" when "1000011001",
      "01010000111100100001001101001011111010011111011000" when "1000011010",
      "01011010111001111000111001110010110110100111111111" when "1000011011",
      "01100100110111111000011101001000010001110100001011" when "1000011100",
      "01101110110110011111111001101011101011111100110110" when "1000011101",
      "01111000110101101111010001111100101110111001001011" when "1000011110",
      "10000010110101100110101000011011001110011111010011" when "1000011111",
      "00001100110110000101111111100111001000100100110111" when "1000100000",
      "00010110110111001101011010000000100100111111101111" when "1000100001",
      "00100000111000111100111010000111110101100110100101" when "1000100010",
      "00101010111011010100100010011101010110010001011100" when "1000100011",
      "00110100111110010100010101100001101100111010011110" when "1000100100",
      "00111111000001111100010101110101101001011110100000" when "1000100101",
      "01001001000110001100100101111010000101111101101010" when "1000100110",
      "01010011001011000101001000010000000110011011111111" when "1000100111",
      "00011101010000100101111111011000111001000010001010" when "1000101000",
      "00100111010110101111001101110101110101111110000000" when "1000101001",
      "00110001011101100000110110001000011111100011001010" when "1000101010",
      "00111011100100111010111010110010100010001011110010" when "1000101011",
      "01000101101100111101011110010101110100011001000101" when "1000101100",
      "01001111110101101000100011010100010110110100000000" when "1000101101",
      "01011001111110111100001100010000010100001101110101" when "1000101110",
      "01100100001000111000011011101100000001100000110110" when "1000101111",
      "00101110010011011101010100001001111101110000111111" when "1000110000",
      "00111000011110101010111000001100110010001100011010" when "1000110001",
      "01000010101010100001001010010111010010001100001010" when "1000110010",
      "01001100110111000000001101001100011011010100110111" when "1000110011",
      "01010111000100001000000011001111010101010111010000" when "1000110100",
      "01100001010001111000101111000011010010010000111010" when "1000110101",
      "01101011100000010010010011001011101110001100110110" when "1000110110",
      "01110101101111010100110010001100001111100100001000" when "1000110111",
      "00111111111111000000001110101000100110111110100101" when "1000111000",
      "01001010001111010100101011000100101111010011010110" when "1000111001",
      "01010100100000010010001010000100101101101001100111" when "1000111010",
      "01011110110001111000101110001100110001011001001010" when "1000111011",
      "01101001000100001000011010000001010100001011000101" when "1000111100",
      "01110011010111000001010000000110111001111010011010" when "1000111101",
      "01111101101010100011010011000010010000110100101011" when "1000111110",
      "10000111111110101110100101011000010001011010101101" when "1000111111",
      "00010010010011100011001001101101111110100001000111" when "1001000000",
      "00011100101001000001000010101000100101010001000010" when "1001000001",
      "00100110111111001000010010101101011101001000110010" when "1001000010",
      "00110001010101111000111100100010000111111100011010" when "1001000011",
      "00111011101101010011000010101100010001110110011010" when "1001000100",
      "01000110000101010110100111110001110001011000011010" when "1001000101",
      "01010000011110000011101110011000100111011011101110" when "1001000110",
      "01011010110111011010011001000110111111010010000010" when "1001000111",
      "00100101010001011010101010100011001110100110000111" when "1001001000",
      "00101111101100000100100101010011110101011100010110" when "1001001001",
      "00111010000111011000001011111111011110010011011111" when "1001001010",
      "01000100100011010101100001001100111110000101010001" when "1001001011",
      "01001110111111111100100111100011010100000111000010" when "1001001100",
      "01011001011101001101100001101001101010001010011100" when "1001001101",
      "01100011111011001000010010000111010100011110000100" when "1001001110",
      "01101110011001101100111011100011110001101110000011" when "1001001111",
      "00111000111000111011100000100110101011000100110110" when "1001010000",
      "01000011011000110100000011110111110100001011110001" when "1001010001",
      "01001101111001010110100111111111001011001011101010" when "1001010010",
      "01011000011010100011001111100100111000101101101000" when "1001010011",
      "01100010111100011001111101010001001111111011100111" when "1001010100",
      "01101101011110111010110011101100101110100001000110" when "1001010101",
      "01111000000010000101110101011111111100101011101111" when "1001010110",
      "10000010100101111011000101010011101101001100000011" when "1001010111",
      "00001101001010011010100101110000111101010110000010" when "1001011000",
      "00010111101111100100011001100000110101000001111000" when "1001011001",
      "00100010010101011000100011001100100110101100100010" when "1001011010",
      "00101100111011110111000101011101101111011000100001" when "1001011011",
      "00110111100011000000000010111101110110101110011011" when "1001011100",
      "01000010001010110011011110010110101110111101101100" when "1001011101",
      "01001100110011010001011010010010010100111101001111" when "1001011110",
      "01010111011100011001111001011010110000001100000101" when "1001011111",
      "00100010000110001100111110011010010010110010000101" when "1001100000",
      "00101100110000101010101011111011011001100000100001" when "1001100001",
      "00110111011011110011000100101000101011110010110101" when "1001100010",
      "01000010000111100110001011001100111011101111010001" when "1001100011",
      "01001100110100000100000010010011000110000111100000" when "1001100100",
      "01010111100001001100101100100110010010011001011001" when "1001100101",
      "01100010001111000000001100110001110010101111100011" when "1001100110",
      "01101100111101011110100101100001000100000010000101" when "1001100111",
      "00110111101100100111111001011111101101110111001110" when "1001101000",
      "01000010011100011100001011011001100010100100000010" when "1001101001",
      "01001101001100111011011101111010011111001101000010" when "1001101010",
      "01010111111110000101110011101110101011100110111011" when "1001101011",
      "01100010101111111011001111100010011010010111001100" when "1001101100",
      "01101101100010011011110100000010001000110100111000" when "1001101101",
      "01111000010101100111100011111010011111001001001000" when "1001101110",
      "10000011001001011110100001111000010000001111111111" when "1001101111",
      "00001101111110000000110000101000011001111000111111" when "1001110000",
      "00011000110011001110010010111000000100100111111001" when "1001110001",
      "00100011101001000111001011010100100011110101010100" when "1001110010",
      "00101110011111101011011100101011010101101111011011" when "1001110011",
      "00111001010110111011001001101010000011011010100111" when "1001110100",
      "01000100001110110110010100111110100000110010001011" when "1001110101",
      "01001111000111011101000001010110101100101001000000" when "1001110110",
      "01011010000000101111010001100000110000101010010000" when "1001110111",
      "00100100111010101101001000001011000001011010000000" when "1001111000",
      "00101111110101010110101000000011111110010110000000" when "1001111001",
      "00111010110000101011110011111010010001110110010001" when "1001111010",
      "01000101101100101100101110011100110001001101110100" when "1001111011",
      "01010000101001011001011010011010011100101011010101" when "1001111100",
      "01011011100110110001111010100010011111011001111000" when "1001111101",
      "01100110100100110110010001100100001111100001100001" when "1001111110",
      "01110001100011100110100010001111001110001000000111" when "1001111111",
      "00111100100011000010101111010011000111010001110101" when "1010000000",
      "01000111100011001010111011011111110010000010000010" when "1010000001",
      "01010010100011111111001001100101010000011011110101" when "1010000010",
      "01011101100101011111011100010011101111100010110001" when "1010000011",
      "01101000100111101011110110011011100111011011100111" when "1010000100",
      "01110011101010100100011010101101011011001100111100" when "1010000101",
      "01111110101110001001001011111001111000111111111000" when "1010000110",
      "10001001110010011010001100110001111010000000110010" when "1010000111",
      "00010100110111010111100000000110100010011111111100" when "1010001000",
      "00011111111101000001001000101001000001110010001111" when "1010001001",
      "00101011000011010111001001001010110010010001110110" when "1010001010",
      "00110110001010011001100100011101011001011110111111" when "1010001011",
      "01000001010010001000011101010010101000000000100001" when "1010001100",
      "01001100011010100011110110011100011001100100101101" when "1010001101",
      "01010111100011101011110010101100110101000001111010" when "1010001110",
      "01100010101101100000010100110110001100010111001111" when "1010001111",
      "00101101111000000001011111101010111100101101010011" when "1010010000",
      "00111001000011001111010101111101101110010110110110" when "1010010001",
      "01000100001111001001111010100001010100110001100001" when "1010010010",
      "01001111011011110001010000001000101110100110100001" when "1010010011",
      "01011010101001000101011001100111000101101011010010" when "1010010100",
      "01100101110111000110011001101111101111000010010000" when "1010010101",
      "01110001000101110100010011010110001010111011100010" when "1010010110",
      "01111100010101001111001001001110000100110101100101" when "1010010111",
      "00000111100101010110111110001011010011011101111010" when "1010011000",
      "00010010110110001011110101000001111000110001110100" when "1010011001",
      "00011110000111101101110000100110000001111111000100" when "1010011010",
      "00101001011001111100110011101100000111100100101001" when "1010011011",
      "00110100101100111001000001001000101101010011010110" when "1010011100",
      "01000000000000100010011011110000100010001110100111" when "1010011101",
      "01001011010100111001000110011000100000101101001001" when "1010011110",
      "01010110101001111101000011110101101110011001101011" when "1010011111",
      "00100001111111101110010110111101011100010011100111" when "1010100000",
      "00101101010110001101000010100101000110101111110011" when "1010100001",
      "00111000101101011001001001100010010101011001001101" when "1010100010",
      "01000100000101010010101110101010111011010001100111" when "1010100011",
      "01001111011101111001110100110100110110110010011001" when "1010100100",
      "01011010110111001110011110110110010001101101000111" when "1010100101",
      "01100110010001010000101111100101100001001100010111" when "1010100110",
      "01110001101100000000101001111001000101110100010111" when "1010100111",
      "00111101000111011110010000100111101011100011110001" when "1010101000",
      "01001000100011101001100110101000001001110100010100" when "1010101001",
      "01010100000000100010101110110001100011011011100011" when "1010101010",
      "01011111011110001001101011111011000110101011100110" when "1010101011",
      "01101010111100011110100000111100001101010011110010" when "1010101100",
      "01110110011011100001010000101100011100100001011011" when "1010101101",
      "10000001111011010001111110000011100101000000100010" when "1010101110",
      "10001101011011110000101011111001100010111100100000" when "1010101111",
      "00011000111100111101011101000110011110000000110101" when "1010110000",
      "00100100011110111000010100100010101001011001111010" when "1010110001",
      "00110000000001100001010101000110100011110101101001" when "1010110010",
      "00111011100100111000100001101010110111100100010000" when "1010110011",
      "01000111001000111101111101001000011010011000111010" when "1010110100",
      "01010010101101110001101010011000001101101010100011" when "1010110101",
      "01011110010011010011101100010011011110010100100011" when "1010110110",
      "01101001111001100100000101110011100100110111011101" when "1010110111",
      "00110101100000100010111001110010000101011001101100" when "1010111000",
      "01000001001000010000001011001000101111101000010100" when "1010111001",
      "01001100110000101011111100110001011110110111101111" when "1010111010",
      "01011000011001110110010001100110011010000100011011" when "1010111011",
      "01100100000011101111001100100001110011110011101000" when "1010111100",
      "01101111101110010110110000011110001010010100001010" when "1010111101",
      "01111011011001101101000000010110000111011111000011" when "1010111110",
      "10000111000101110001111111000100100000111000010101" when "1010111111",
      "00010010110010100101101111100100010111101111110001" when "1011000000",
      "00011110100000001000010100110000111001000001100001" when "1011000001",
      "00101010001110011001110001100101011101010110111100" when "1011000010",
      "00110101111101011010001000111101101001000111010101" when "1011000011",
      "01000001101101001001011101110101001100011000100100" when "1011000100",
      "01001101011101100111110011001000000010111111111100" when "1011000101",
      "01011001001110110101001011110010010100100010110101" when "1011000110",
      "01100101000000110001101010110000010100010111011101" when "1011000111",
      "00110000110011011101010010111110100001100101101001" when "1011001000",
      "00111100100110111000000111011001100111000111011111" when "1011001001",
      "01001000011011000010001010111110011011101010001011" when "1011001010",
      "01010100001111111011100000101010000001101110101001" when "1011001011",
      "01100000000101100100001011011001100111101010011000" when "1011001100",
      "01101011111011111100001110001010100111101000001000" when "1011001101",
      "01110111110011000011101011111010100111101000101010" when "1011001110",
      "10000011101010111010100111100111011001100011011101" when "1011001111",
      "00001111100011100001000100001110111011000111100000" when "1011010000",
      "00011011011100110111000100101111010101111100000001" when "1011010001",
      "00100111010110111100101100000110111111100001001101" when "1011010010",
      "00110011010001110001111101010100011001010000111101" when "1011010011",
      "00111111001101010110111011010110010000011111101001" when "1011010100",
      "01001011001001101011101001001011011110011100110100" when "1011010101",
      "01010111000110110000001001110011001000010100000001" when "1011010110",
      "01100011000100100100100000001100011111001101011101" when "1011010111",
      "00101111000011001000101111010111000000001110110010" when "1011011000",
      "00111011000010011100111010010010010100011011111000" when "1011011001",
      "01000111000010100001000011111110010000110111100000" when "1011011010",
      "01010011000011010101001111011010110110100100001011" when "1011011011",
      "01011111000100111001011111101000010010100100110010" when "1011011100",
      "01101011000111001101110111100110111101111101011110" when "1011011101",
      "01110111001010010010011010010111011101110100010010" when "1011011110",
      "10000011001110000111001010111010100011010001111110" when "1011011111",
      "00001111010010101100001100010001001011100010101111" when "1011100000",
      "00011011011000000001100001011100011111110110111111" when "1011100001",
      "00100111011110000111001101011101110101100100000101" when "1011100010",
      "00110011100100111101010011010110101110000101000100" when "1011100011",
      "00111111101100100011110110001000110110111011100000" when "1011100100",
      "01001011110100111010111000110110001001110000001001" when "1011100101",
      "01010111111110000010011110100000101100010011101101" when "1011100110",
      "01100100000111111010101010001010110000011111101101" when "1011100111",
      "00110000010010100011011110110110110100010111000101" when "1011101000",
      "00111100011101111100111111100111100010000111000111" when "1011101001",
      "01001000101010000111001111011111110000001000000001" when "1011101010",
      "01010100110111000010010001100010100000111101110110" when "1011101011",
      "01100001000100101110001000110011000011011001001010" when "1011101100",
      "01101101010011001010111000010100110010010111110110" when "1011101101",
      "01111001100010011000100011001011010101000101110111" when "1011101110",
      "10000101110010010111001100011010011110111101111101" when "1011101111",
      "00010010000011000110110111000110001111101010100010" when "1011110000",
      "00011110010100100111100110010010110011000110010011" when "1011110001",
      "00101010100110111001011101000100100001011101001001" when "1011110010",
      "00110110111001111100011110011111111111001100110011" when "1011110011",
      "01000011001101110000101101101001111101000101101101" when "1011110100",
      "01001111100010010110001101100111011000001011101101" when "1011110101",
      "01011011110111101101000001011101011001110110110110" when "1011110110",
      "01101000001101110101001100010001010111110100001011" when "1011110111",
      "00110100100100101110110001001000110100000110011101" when "1011111000",
      "01000000111100011001110011001001011101000110111100" when "1011111001",
      "01001101010100110110010101011001001101100110001111" when "1011111010",
      "01011001101110000100011010111110001100101100111100" when "1011111011",
      "01100110001000000100000110111110101101111100100010" when "1011111100",
      "01110010100010110101011100100001010001010000000011" when "1011111101",
      "01111110111110011000011110101100100010111100111110" when "1011111110",
      "10001011011010101101010000100111011011110011111001" when "1011111111",
      "00010111110111110011110101011001000001000001010111" when "1100000000",
      "00100100010101101100010000001000100100001110101001" when "1100000001",
      "00110000110100010110100011111101100011100010011110" when "1100000010",
      "00111101010011110010110011111111101001100001111000" when "1100000011",
      "01001001110100000001000011010110101101010000111100" when "1100000100",
      "01010110010101000001010101001010110010010011100011" when "1100000101",
      "01100010110110110011101100100100001000101110010000" when "1100000110",
      "01101111011001011000001100101011001101000110111011" when "1100000111",
      "00111011111100101110111000101000101000100101101100" when "1100001000",
      "01001000100000110111110011100101010000110101100110" when "1100001001",
      "01010101000101110011000000101010001000000101011100" when "1100001010",
      "01100001101011100000100011000000011101001000100011" when "1100001011",
      "01101110010010000000011101110001101011010111100110" when "1100001100",
      "01111010111001010010110100000111011010110001010100" when "1100001101",
      "10000111100001010111101001001011011111111011011000" when "1100001110",
      "10010100001010001111000000000111111100000011000111" when "1100001111",
      "00100000110011111000111100000110111100111110010100" when "1100010000",
      "00101101011110010101100000010010111101001100000011" when "1100010001",
      "00111010001001100100101111110110100011110101011011" when "1100010010",
      "01000110110101100110101101111100100100101110011001" when "1100010011",
      "01010011100010011011011101110000000000010110100100" when "1100010100",
      "01100000010000000011000010011100000011111001111011" when "1100010101",
      "01101100111110011101011111001100001001010001101111" when "1100010110",
      "01111001101101101010110111001011110111000101010000" when "1100010111",
      "00000110011101101011001101100111000000101010100010" when "1100011000",
      "00010011001110011110100101101001100110000111001111" when "1100011001",
      "00100000000000000101000010011111110100010001011110" when "1100011010",
      "00101100110010011110100111010110000100110000011111" when "1100011011",
      "00111001100101101011010111011000111101111101100100" when "1100011100",
      "01000110011001101011010101110101010011000100110011" when "1100011101",
      "01010011001110011110100101111000000100000101110111" when "1100011110",
      "01100000000100000101001010101110011101110100110100" when "1100011111",
      "00101100111010011111000111100101111001111010111101" when "1100100000",
      "00111001110001101100011111101011111110110111100100" when "1100100001",
      "01000110101001101101010110001110100000000000101111" when "1100100010",
      "01010011100010100001101110011011011101100100001010" when "1100100011",
      "01100000011100001001101011100001000100100111111101" when "1100100100",
      "01101101010110100101010000101101101111001011011101" when "1100100101",
      "01111010010001110100100001010000000100001000000011" when "1100100110",
      "10000111001101110111100000010110110111010001111011" when "1100100111",
      "00010100001010101110010001010001001001011000111100" when "1100101000",
      "00100001001000011000110111001110001000001001010111" when "1100101001",
      "00101110000110110111010101011101001110001100110001" when "1100101010",
      "00111011000110001001101111001110000011001010110001" when "1100101011",
      "01001000000110010000000111110000011011101001111001" when "1100101100",
      "01010101000111001010100010010100011001010000010101" when "1100101101",
      "01100010001000111001000010001010001010100100110010" when "1100101110",
      "01101111001011011011101010100010001011001111010010" when "1100101111",
      "00111100001110110010011110101101000011111010000000" when "1100110000",
      "01001001010010111101100001111011101010010010000011" when "1100110001",
      "01010110010111111100110111011111000001001000010011" when "1100110010",
      "01100011011101110000100010101000011000010010001100" when "1100110011",
      "01110000100100011000100110101001001100101010100110" when "1100110100",
      "01111101101011110101000110110011001000010010100101" when "1100110101",
      "10001010110100000110000110011000000010010010010000" when "1100110110",
      "10010111111101001011101000101001111110111001100101" when "1100110111",
      "00100101000111000101110000111011001111100001001100" when "1100111000",
      "00110010010001110100100010011110010010101011001111" when "1100111001",
      "00111111011101011000000000100101110100000100001001" when "1100111010",
      "01001100101001110000001110100100101100100011100011" when "1100111011",
      "01011001110110111101001111101110000010001100111111" when "1100111100",
      "01100111000100111111000111010101001000010000110100" when "1100111101",
      "01110100010011110101111000101101011111001101000010" when "1100111110",
      "10000001100011100001100111001010110100101110000001" when "1100111111",
      "00001110110100000010010110000001000011101111011110" when "1101000000",
      "00011100000101011000001000100100010100011101001011" when "1101000001",
      "00101001010111100011000010001000111100010011110101" when "1101000010",
      "00110110101010100011000110000011011110000001111010" when "1101000011",
      "01000011111110011000010111101000101001101000011101" when "1101000100",
      "01010001010011000010111010001101011100011011111011" when "1101000101",
      "01011110101000100010110001000111000001000101000010" when "1101000110",
      "01101011111110110111111111101010101111100001100101" when "1101000111",
      "00111001010110000010101001001110001101000101010010" when "1101001000",
      "01000110101110000010110001000111001100011010100101" when "1101001001",
      "01010100000110111000011010101011101101100011100010" when "1101001010",
      "01100001100000100011101001010001111101111010100101" when "1101001011",
      "01101110111011000100100000010000011000010011011110" when "1101001100",
      "01111100010110011011000010111101100100111011111111" when "1101001101",
      "10001001110010100111010100110000011001011100111010" when "1101001110",
      "10010111001111101001011000111111111000111010101110" when "1101001111",
      "00100100101101100001010011000011010011110110100101" when "1101010000",
      "00110010001100001111000110010010001000001111000100" when "1101010001",
      "00111111101011110010110110000100000001100001000010" when "1101010010",
      "01001101001100001100100101110000111000101000100010" when "1101010011",
      "01011010101101011100011000110000110100000001100010" when "1101010100",
      "01101000001111100010010010011100000111101000110111" when "1101010101",
      "01110101110010011110010110001011010100111101000001" when "1101010110",
      "10000011010110010000100111010111001010111110111111" when "1101010111",
      "00010000111010111001001001011000100110010011001010" when "1101011000",
      "00011110100000010111111111101000110001000010000101" when "1101011001",
      "00101100000110101101001101100001000010111001011011" when "1101011010",
      "00111001101101111000110110011011000001001100101100" when "1101011011",
      "01000111010101111010111101110000011110110110001110" when "1101011100",
      "01010100111110110011100110111011011100010111111000" when "1101011101",
      "01100010101000100010110101010110000111111100000011" when "1101011110",
      "01110000010011001000101100011010111101010110011001" when "1101011111",
      "00111101111110100101001111100100100110000100110001" when "1101100000",
      "01001011101010111000100010001101111001010000000010" when "1101100001",
      "01011001011000000010100111110001111011101100111010" when "1101100010",
      "01100111000110000011100011101011111111111100110111" when "1101100011",
      "01110100110100111011011001010111100110001110111011" when "1101100100",
      "10000010100100101010001100010000011100100000101000" when "1101100101",
      "10010000010101001111111111110010011110011110101110" when "1101100110",
      "10011110000110101100110111011001110101100110001101" when "1101100111",
      "00101011111001000000110110100010111001000101000000" when "1101101000",
      "00111001101100001100000000101010001101111011000001" when "1101101001",
      "01000111100000001110011001001100100110111010110101" when "1101101010",
      "01010101010101001000000011100111000100101010101001" when "1101101011",
      "01100011001010111001000011010110110101100101001000" when "1101101100",
      "01110001000001100001011011111001010101111010010100" when "1101101101",
      "01111110111001000001010000101100001111110000011001" when "1101101110",
      "10001100110001011000100101001101011011000100101001" when "1101101111",
      "00011010101010100111011100111010111101101100010000" when "1101110000",
      "00101000100100101101111011010011001011010101001111" when "1101110001",
      "00110110011111101100000011110100100101100111010000" when "1101110010",
      "01000100011011100001111001111101111100000100100001" when "1101110011",
      "01010010011000001111100001001110001100001010101000" when "1101110100",
      "01100000010101110100111101000100100001010011011110" when "1101110101",
      "01101110010100010010010001000000010100110110000101" when "1101110110",
      "01111100010011100111100000100001001110000111100001" when "1101110111",
      "00001010010011110100101111000111000010011011101110" when "1101111000",
      "00011000010100111010000000010001110101000110011100" when "1101111001",
      "00100110010110110111010111100001110111011100000001" when "1101111010",
      "00110100011001101100111000010111101000110010010110" when "1101111011",
      "01000010011101011010100110010011110110100001101100" when "1101111100",
      "01010000100010000000100100110111011100000101101001" when "1101111101",
      "01011110100111011110110111100011100010111101111001" when "1101111110",
      "01101100101101110101100001111001100010101111001100" when "1101111111",
      "00111010110101000100100111011011000001000100001100" when "1110000000",
      "01001000111101001100001011101001110001101110010111" when "1110000001",
      "01010111000110001100010010000111110110100110110100" when "1110000010",
      "01100101010000000100111110010111011111101111010001" when "1110000011",
      "01110011011010110110010011111011001011010010110101" when "1110000100",
      "10000001100110100000010110010101100101100110111110" when "1110000101",
      "10001111110011000011001001001001101001001100011000" when "1110000110",
      "10011110000000011110101111111010011110101111110100" when "1110000111",
      "00101100001110110011001110001011011101001011000100" when "1110001000",
      "00111010011110000000100111100000001001100101110000" when "1110001001",
      "01001000101110000110111111011100010111010110010010" when "1110001010",
      "01010110111111000110011001100100001000000010101110" when "1110001011",
      "01100101010000111110111001011011101011100001101011" when "1110001100",
      "01110011100011110000100010100111011111111011001011" when "1110001101",
      "10000001110111011011011000101100010001101001100110" when "1110001110",
      "10010000001011111111011111001110111011011010100010" when "1110001111",
      "00011110100001011100111001110100100110001111101101" when "1110010000",
      "00101100110111110011101100000010101001011111110100" when "1110010001",
      "00111011001111000011111001011110101010110111100000" when "1110010010",
      "01001001100111001101100101101110011110011010001101" when "1110010011",
      "01011000000000010000110100011000000110100011000100" when "1110010100",
      "01100110011010001101101001000001110100000101110011" when "1110010101",
      "01110100110101000100000111010010000110001111101010" when "1110010110",
      "10000011010000110100010010101111101010101000010010" when "1110010111",
      "00010001101101011110001111000001011101010010100111" when "1110011000",
      "00100000001011000001111111101110101000101101110010" when "1110011001",
      "00101110101001011111101000011110100101110110000011" when "1110011010",
      "00111101001000110111001100111000111100000101101100" when "1110011011",
      "01001011101001001000110000100101100001010101110111" when "1110011100",
      "01011010001010010100010111001100011001111111100101" when "1110011101",
      "01101000101100011010000100010101111000111100100100" when "1110011110",
      "01110111001111011001111011101010011111101000001100" when "1110011111",
      "00000101110011010100000000110010111110000000010110" when "1110100000",
      "00010100011000001000010111011000010010100110011001" when "1110100001",
      "00100010111101110111000011000011101010100000000011" when "1110100010",
      "00110001100100100000000111011110100001011000010101" when "1110100011",
      "01000000001100000011101000010010100001100000011010" when "1110100100",
      "01001110110100100001101001001001100011110000100100" when "1110100101",
      "01011101011101111010001101101101101111101001000100" when "1110100110",
      "01101100001000001101011001101001011011010011001011" when "1110100111",
      "00111010110011011011010000100111001011100001111010" when "1110101000",
      "01001001011111100011110110010001110011110011000110" when "1110101001",
      "01011000001100100111001110010100010110010000010000" when "1110101010",
      "01100110111010100101011100011010000011101111011100" when "1110101011",
      "01110101101001011110100100001110011011110100010000" when "1110101100",
      "10000100011001010010101001011101001100110000110000" when "1110101101",
      "10010011001010000001101111110010010011100110010011" when "1110101110",
      "10100001111011101011111010111001111100000110100100" when "1110101111",
      "00110000101110010001001110100000100000110100011001" when "1110110000",
      "00111111100001110001101110010010101011000100110001" when "1110110001",
      "01001110010110001101011101111101010010111111101110" when "1110110010",
      "01011101001011100100100001001101011111100001001110" when "1110110011",
      "01101100000001110110111011110000100110011010001100" when "1110110100",
      "01111010111001000100110001010100001100010001010101" when "1110110101",
      "10001001110001001110000101100110000100100100000110" when "1110110110",
      "10011000101010010010111100010100010001100111101010" when "1110110111",
      "00100111100100010011011001001101000100101001110000" when "1110111000",
      "00110110011111001111011111111110111101110001101100" when "1110111001",
      "01000101011011000111010100011000101100000001001111" when "1110111010",
      "01010100010111111010111010001001001101010101100101" when "1110111011",
      "01100011010101101010010100111111101110101000001110" when "1110111100",
      "01110010010100010101101000101011101011101111111110" when "1110111101",
      "10000001010011111100111000111100101111100001110100" when "1110111110",
      "10010000010100100000001001100010110011110001111010" when "1110111111",
      "00011111010101111111011110001110000001010100011110" when "1111000000",
      "00101110011000011010111010101110101111111110110000" when "1111000001",
      "00111101011011110010100010110101100110100111111110" when "1111000010",
      "01001100100000000110011010010011011011001010001101" when "1111000011",
      "01011011100101010110100100111001010010100011011010" when "1111000100",
      "01101010101011100011000110011000100000110110010100" when "1111000101",
      "01111001110010101100000010100010101001001011011000" when "1111000110",
      "10001000111010110001011101001001011101110001101101" when "1111000111",
      "00011000000011110011011001111111000000000000000011" when "1111001000",
      "00100111001101110001111100110101100000010101101010" when "1111001001",
      "00110110011000101101001001011111011110011011010111" when "1111001010",
      "01000101100100100101000011101111101001000100011000" when "1111001011",
      "01010100110001011001101111011000111110001111011000" when "1111001100",
      "01100011111111001011010000001110101011000111010100" when "1111001101",
      "01110011001101111001101010000100001100000100100000" when "1111001110",
      "10000010011101100101000000101101001100101101011110" when "1111001111",
      "00010001101110001101010111111101100111110111111110" when "1111010000",
      "00100000111111110010110011101001100111101001111000" when "1111010001",
      "00110000010010010101010111100101100101011010001101" when "1111010010",
      "00111111100101110101000111100110001001110010000001" when "1111010011",
      "01001110111010010010000111100000001100101101011000" when "1111010100",
      "01011110001111101100011011001000110101011100011000" when "1111010101",
      "01101101100110000100000110010101011010100011111110" when "1111010110",
      "01111100111101011001001100111011100001111111000100" when "1111010111",
      "00001100010101101011110010110001000000111111011000" when "1111011000",
      "00011011101110111011111011101011111100001110011100" when "1111011001",
      "00101011001001001001101011100010100111101110100100" when "1111011010",
      "00111010100100010101000110001011100110111011110011" when "1111011011",
      "01001010000000011110001111011101101100101100111001" when "1111011100",
      "01011001011101100101001011001111111011010100001110" when "1111011101",
      "01101000111011101001111101011001100100100000110110" when "1111011110",
      "01111000011010101100101001110010001001011111010111" when "1111011111",
      "00000111111010101101010100010001011010111010111101" when "1111100000",
      "00010111011011101100000000101111011000111110010100" when "1111100001",
      "00100110111101101000110011000100010011010100101001" when "1111100010",
      "00110110100000100011101111001000101001001010101000" when "1111100011",
      "01000110000100011100111000110101001001001111010101" when "1111100100",
      "01010101101001010100010100000010110001110101010010" when "1111100101",
      "01100101001111001010000100101010110000110011010110" when "1111100110",
      "01110100110101111110001110100110100011100101110010" when "1111100111",
      "00000100011101110000110101101111110111001111001001" when "1111101000",
      "00010100000110100001111110000000101000011001010010" when "1111101001",
      "00100011110000010001101011010011000011010110011000" when "1111101010",
      "00110011011011000000000001100001100100000001110100" when "1111101011",
      "01000011000110101101000100100110110110000001001111" when "1111101100",
      "01010010110011011000111000011101110100100101011111" when "1111101101",
      "01100010100001000011100001000001101010101011100111" when "1111101110",
      "01110010001111101101000010001101110010111101110111" when "1111101111",
      "00000001111111010101011111111101110111110100100101" when "1111110000",
      "00010001101111111100111110001101110011010111010011" when "1111110001",
      "00100001100001100011100000111001101111011101101010" when "1111110010",
      "00110001010100001001001011111110000101110000011011" when "1111110011",
      "01000001000111101110000011010111011111101010011100" when "1111110100",
      "01010000111100010010001011000010110110011001101001" when "1111110101",
      "01100000110001110101100110111101010011000000000001" when "1111110110",
      "01110000101000011000011011000100001110010100101001" when "1111110111",
      "00000000011111111010101011010101010001000100101000" when "1111111000",
      "00010000011000011100011011101110010011110100000110" when "1111111001",
      "00100000010001111101110000001101011110111111010001" when "1111111010",
      "00110000001100011110101100110001001010111011010100" when "1111111011",
      "01000000000111111111010101010111111111110111011110" when "1111111100",
      "01010000000100011111101110000000110101111101111110" when "1111111101",
      "01100000000001111111111010101010110101010101000100" when "1111111110",
      "01110000000000011111111111010101010101111111111111" when "1111111111",
      "--------------------------------------------------" when others;
   Y1_c19 <= Y0_c19; -- for the possible blockram register
   Y <= Y1_c19;
end architecture;

--------------------------------------------------------------------------------
--                      compressedTable_Freq300_uid1527
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Luc Forget, Maxime Christ (2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq300_uid1527 is
    port (clk, ce_20 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of compressedTable_Freq300_uid1527 is
   component compressedTable_Freq300_uid1527_subsampling_Freq300_uid1529 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(8 downto 0)   );
   end component;

   component compressedTable_Freq300_uid1527_diff_Freq300_uid1532 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(49 downto 0)   );
   end component;

signal X_subsampling_c19 :  std_logic_vector(6 downto 0);
signal Y_subsampling_c19, Y_subsampling_c20 :  std_logic_vector(8 downto 0);
signal Y_subsampling_copy1530_c19 :  std_logic_vector(8 downto 0);
signal Y_diff_c19, Y_diff_c20 :  std_logic_vector(49 downto 0);
signal fullOut_topbits_c20 :  std_logic_vector(8 downto 0);
signal fullOut_c20 :  std_logic_vector(56 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               Y_subsampling_c20 <= Y_subsampling_c19;
               Y_diff_c20 <= Y_diff_c19;
            end if;
         end if;
      end process;
   X_subsampling_c19 <= X(9 downto 3);
   compressedTable_Freq300_uid1527_subsampling: compressedTable_Freq300_uid1527_subsampling_Freq300_uid1529
      port map ( X => X_subsampling_c19,
                 Y => Y_subsampling_copy1530_c19);
   Y_subsampling_c19 <= Y_subsampling_copy1530_c19; -- output copy to hold a pipeline register if needed
   compressedTable_Freq300_uid1527_diff: compressedTable_Freq300_uid1527_diff_Freq300_uid1532
      port map ( clk  => clk,
                 X => X,
                 Y => Y_diff_c19);
   fullOut_topbits_c20 <= Y_subsampling_c20 + ("0000000"& (Y_diff_c20(49 downto 48)));
   fullOut_c20 <= fullOut_topbits_c20 & (Y_diff_c20(47 downto 0));
   Y <= fullOut_c20;
end architecture;

--------------------------------------------------------------------------------
--                     FixFunctionByTable_Freq300_uid1525
-- Evaluator for exp(x*1b-1) on [-1,1) for lsbIn=-9 (wIn=10), msbout=0, lsbOut=-56 (wOut=57). Out interval: [0.606531; 1.64711]. Output is unsigned

-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq300_uid1525 is
    port (clk, ce_20 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq300_uid1525 is
   component compressedTable_Freq300_uid1527 is
      port ( clk, ce_20 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(56 downto 0)   );
   end component;

begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
            end if;
         end if;
      end process;
   compressedTable: compressedTable_Freq300_uid1527
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 X => X,
                 Y => Y);
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid1544
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid1544 is
    port (clk, ce_20 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid1544 is
signal Mfull_c19, Mfull_c20 :  std_logic_vector(40 downto 0);
signal M_c20 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               Mfull_c20 <= Mfull_c19;
            end if;
         end if;
      end process;
   Mfull_c19 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c20 <= Mfull_c20(40 downto 0);
   R <= M_c20;
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1546
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1546 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1546 is
   component MultTable_Freq300_uid1548 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1549_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1548
      port map ( X => Xtable_c19,
                 Y => Y1_copy1549_c19);
   Y1_c19 <= Y1_copy1549_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1551
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1551 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1551 is
   component MultTable_Freq300_uid1553 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1554_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1553
      port map ( X => Xtable_c19,
                 Y => Y1_copy1554_c19);
   Y1_c19 <= Y1_copy1554_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1556
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1556 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1556 is
   component MultTable_Freq300_uid1558 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1559_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1558
      port map ( X => Xtable_c19,
                 Y => Y1_copy1559_c19);
   Y1_c19 <= Y1_copy1559_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1561
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1561 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1561 is
   component MultTable_Freq300_uid1563 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1564_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1563
      port map ( X => Xtable_c19,
                 Y => Y1_copy1564_c19);
   Y1_c19 <= Y1_copy1564_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1566
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1566 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1566 is
   component MultTable_Freq300_uid1568 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1569_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1568
      port map ( X => Xtable_c19,
                 Y => Y1_copy1569_c19);
   Y1_c19 <= Y1_copy1569_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1571
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1571 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1571 is
   component MultTable_Freq300_uid1573 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1574_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1573
      port map ( X => Xtable_c19,
                 Y => Y1_copy1574_c19);
   Y1_c19 <= Y1_copy1574_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1576
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1576 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1576 is
   component MultTable_Freq300_uid1578 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1579_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1578
      port map ( X => Xtable_c19,
                 Y => Y1_copy1579_c19);
   Y1_c19 <= Y1_copy1579_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1581
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1581 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1581 is
   component MultTable_Freq300_uid1583 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1584_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1583
      port map ( X => Xtable_c19,
                 Y => Y1_copy1584_c19);
   Y1_c19 <= Y1_copy1584_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1586
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1586 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1586 is
   component MultTable_Freq300_uid1588 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1589_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1588
      port map ( X => Xtable_c19,
                 Y => Y1_copy1589_c19);
   Y1_c19 <= Y1_copy1589_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1591
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1591 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1591 is
   component MultTable_Freq300_uid1593 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1594_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1593
      port map ( X => Xtable_c19,
                 Y => Y1_copy1594_c19);
   Y1_c19 <= Y1_copy1594_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1596
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1596 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1596 is
   component MultTable_Freq300_uid1598 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1599_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1598
      port map ( X => Xtable_c19,
                 Y => Y1_copy1599_c19);
   Y1_c19 <= Y1_copy1599_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1601
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1601 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1601 is
   component MultTable_Freq300_uid1603 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1604_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1603
      port map ( X => Xtable_c19,
                 Y => Y1_copy1604_c19);
   Y1_c19 <= Y1_copy1604_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1606
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1606 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1606 is
   component MultTable_Freq300_uid1608 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1609_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1608
      port map ( X => Xtable_c19,
                 Y => Y1_copy1609_c19);
   Y1_c19 <= Y1_copy1609_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1611
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1611 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1611 is
   component MultTable_Freq300_uid1613 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1614_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1613
      port map ( X => Xtable_c19,
                 Y => Y1_copy1614_c19);
   Y1_c19 <= Y1_copy1614_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1616
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1616 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1616 is
   component MultTable_Freq300_uid1618 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1619_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1618
      port map ( X => Xtable_c19,
                 Y => Y1_copy1619_c19);
   Y1_c19 <= Y1_copy1619_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1621
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1621 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1621 is
   component MultTable_Freq300_uid1623 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1624_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1623
      port map ( X => Xtable_c19,
                 Y => Y1_copy1624_c19);
   Y1_c19 <= Y1_copy1624_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1626
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1626 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1626 is
   component MultTable_Freq300_uid1628 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1629_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1628
      port map ( X => Xtable_c19,
                 Y => Y1_copy1629_c19);
   Y1_c19 <= Y1_copy1629_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1631
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1631 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1631 is
   component MultTable_Freq300_uid1633 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1634_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1633
      port map ( X => Xtable_c19,
                 Y => Y1_copy1634_c19);
   Y1_c19 <= Y1_copy1634_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1636
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1636 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1636 is
   component MultTable_Freq300_uid1638 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1639_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1638
      port map ( X => Xtable_c19,
                 Y => Y1_copy1639_c19);
   Y1_c19 <= Y1_copy1639_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1641
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1641 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1641 is
   component MultTable_Freq300_uid1643 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1644_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1643
      port map ( X => Xtable_c19,
                 Y => Y1_copy1644_c19);
   Y1_c19 <= Y1_copy1644_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1646
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1646 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1646 is
   component MultTable_Freq300_uid1648 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1649_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1648
      port map ( X => Xtable_c19,
                 Y => Y1_copy1649_c19);
   Y1_c19 <= Y1_copy1649_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1651
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1651 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1651 is
   component MultTable_Freq300_uid1653 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1654_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1653
      port map ( X => Xtable_c19,
                 Y => Y1_copy1654_c19);
   Y1_c19 <= Y1_copy1654_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1656
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1656 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1656 is
   component MultTable_Freq300_uid1658 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1659_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1658
      port map ( X => Xtable_c19,
                 Y => Y1_copy1659_c19);
   Y1_c19 <= Y1_copy1659_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1661
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1661 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1661 is
   component MultTable_Freq300_uid1663 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1664_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1663
      port map ( X => Xtable_c19,
                 Y => Y1_copy1664_c19);
   Y1_c19 <= Y1_copy1664_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1666
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1666 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1666 is
   component MultTable_Freq300_uid1668 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1669_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1668
      port map ( X => Xtable_c19,
                 Y => Y1_copy1669_c19);
   Y1_c19 <= Y1_copy1669_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1671
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1671 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1671 is
   component MultTable_Freq300_uid1673 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1674_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1673
      port map ( X => Xtable_c19,
                 Y => Y1_copy1674_c19);
   Y1_c19 <= Y1_copy1674_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1676
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1676 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1676 is
   component MultTable_Freq300_uid1678 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1679_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1678
      port map ( X => Xtable_c19,
                 Y => Y1_copy1679_c19);
   Y1_c19 <= Y1_copy1679_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1681
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1681 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1681 is
   component MultTable_Freq300_uid1683 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1684_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1683
      port map ( X => Xtable_c19,
                 Y => Y1_copy1684_c19);
   Y1_c19 <= Y1_copy1684_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1686
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1686 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1686 is
   component MultTable_Freq300_uid1688 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1689_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1688
      port map ( X => Xtable_c19,
                 Y => Y1_copy1689_c19);
   Y1_c19 <= Y1_copy1689_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1691
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1691 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1691 is
   component MultTable_Freq300_uid1693 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1694_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1693
      port map ( X => Xtable_c19,
                 Y => Y1_copy1694_c19);
   Y1_c19 <= Y1_copy1694_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1696
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1696 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1696 is
   component MultTable_Freq300_uid1698 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1699_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1698
      port map ( X => Xtable_c19,
                 Y => Y1_copy1699_c19);
   Y1_c19 <= Y1_copy1699_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1701
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1701 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1701 is
   component MultTable_Freq300_uid1703 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1704_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1703
      port map ( X => Xtable_c19,
                 Y => Y1_copy1704_c19);
   Y1_c19 <= Y1_copy1704_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1706
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1706 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1706 is
   component MultTable_Freq300_uid1708 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1709_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1708
      port map ( X => Xtable_c19,
                 Y => Y1_copy1709_c19);
   Y1_c19 <= Y1_copy1709_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_2_signedx2_Freq300_uid1711
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid1711 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid1711 is
   component MultTable_Freq300_uid1713 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(3 downto 0);
signal Y1_c19 :  std_logic_vector(3 downto 0);
signal Y1_copy1714_c19 :  std_logic_vector(3 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1713
      port map ( X => Xtable_c19,
                 Y => Y1_copy1714_c19);
   Y1_c19 <= Y1_copy1714_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1716
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1716 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1716 is
   component MultTable_Freq300_uid1718 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1719_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1718
      port map ( X => Xtable_c19,
                 Y => Y1_copy1719_c19);
   Y1_c19 <= Y1_copy1719_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1721
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1721 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1721 is
   component MultTable_Freq300_uid1723 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1724_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1723
      port map ( X => Xtable_c19,
                 Y => Y1_copy1724_c19);
   Y1_c19 <= Y1_copy1724_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_1x1_signed_Freq300_uid1726
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_signed_Freq300_uid1726 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_signed_Freq300_uid1726 is
signal replicated_c19 :  std_logic_vector(0 downto 0);
signal prod_c19 :  std_logic_vector(0 downto 0);
begin
   replicated_c19 <= (0 downto 0 => X(0));
   prod_c19 <= Y and replicated_c19;
   R <= prod_c19;
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid1728
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid1728 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid1728 is
   component MultTable_Freq300_uid1730 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1731_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1730
      port map ( X => Xtable_c19,
                 Y => Y1_copy1731_c19);
   Y1_c19 <= Y1_copy1731_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid1733
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid1733 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid1733 is
   component MultTable_Freq300_uid1735 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1736_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1735
      port map ( X => Xtable_c19,
                 Y => Y1_copy1736_c19);
   Y1_c19 <= Y1_copy1736_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid1738
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid1738 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid1738 is
   component MultTable_Freq300_uid1740 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1741_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1740
      port map ( X => Xtable_c19,
                 Y => Y1_copy1741_c19);
   Y1_c19 <= Y1_copy1741_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid1743
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid1743 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid1743 is
   component MultTable_Freq300_uid1745 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1746_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1745
      port map ( X => Xtable_c19,
                 Y => Y1_copy1746_c19);
   Y1_c19 <= Y1_copy1746_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--             IntMultiplierLUT_4_signedx1_signed_Freq300_uid1748
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4_signedx1_signed_Freq300_uid1748 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4_signedx1_signed_Freq300_uid1748 is
   component MultTable_Freq300_uid1750 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1751_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1750
      port map ( X => Xtable_c19,
                 Y => Y1_copy1751_c19);
   Y1_c19 <= Y1_copy1751_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid1753
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid1753 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid1753 is
   component MultTable_Freq300_uid1755 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c19 :  std_logic_vector(4 downto 0);
signal Y1_c19 :  std_logic_vector(4 downto 0);
signal Y1_copy1756_c19 :  std_logic_vector(4 downto 0);
begin
Xtable_c19 <= Y & X;
   R <= Y1_c19;
   TableMult: MultTable_Freq300_uid1755
      port map ( X => Xtable_c19,
                 Y => Y1_copy1756_c19);
   Y1_c19 <= Y1_copy1756_c19; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_Freq300_uid2009
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_Freq300_uid2009 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_Freq300_uid2009 is
signal Rtmp_c21 :  std_logic_vector(32 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19, Cin_c20, Cin_c21 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               Cin_c19 <= Cin_c18;
            end if;
            if ce_20 = '1' then
               Cin_c20 <= Cin_c19;
            end if;
            if ce_21 = '1' then
               Cin_c21 <= Cin_c20;
            end if;
         end if;
      end process;
   Rtmp_c21 <= X + Y + Cin_c21;
   R <= Rtmp_c21;
end architecture;

--------------------------------------------------------------------------------
--   FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid1541
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan, 2012-2014, 2024
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y A
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid1541 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(24 downto 0);
          Y : in  std_logic_vector(24 downto 0);
          A : in  std_logic_vector(32 downto 0);
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid1541 is
   component DSPBlock_17x24_Freq300_uid1544 is
      port ( clk, ce_20 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1546 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1551 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1556 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1561 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1566 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1571 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1576 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1581 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1586 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1591 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1596 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1601 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1606 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1611 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1616 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1621 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1626 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1631 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1636 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1641 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1646 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1651 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1656 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1661 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1666 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1671 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1676 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1681 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1686 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1691 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1696 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1701 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1706 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid1711 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1716 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1721 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_signed_Freq300_uid1726 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid1728 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid1733 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid1738 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid1743 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4_signedx1_signed_Freq300_uid1748 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid1753 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid1759 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid1763 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid1767 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid1775 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid1809 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_33_Freq300_uid2009 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal XX_c19 :  signed(0+24 downto 0);
signal YY_c19 :  signed(-17+41 downto 0);
signal AA_c19 :  signed(-9+41 downto 0);
signal tile_0_X_c19 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c19 :  std_logic_vector(23 downto 0);
signal tile_0_output_c20 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c20 :  unsigned(40-0 downto 0);
signal bh1542_wm65_0_c20, bh1542_wm65_0_c21 :  std_logic;
signal bh1542_wm64_0_c20, bh1542_wm64_0_c21 :  std_logic;
signal bh1542_wm63_0_c20, bh1542_wm63_0_c21 :  std_logic;
signal bh1542_wm62_0_c20, bh1542_wm62_0_c21 :  std_logic;
signal bh1542_wm61_0_c20, bh1542_wm61_0_c21 :  std_logic;
signal bh1542_wm60_0_c20, bh1542_wm60_0_c21 :  std_logic;
signal bh1542_wm59_0_c20, bh1542_wm59_0_c21 :  std_logic;
signal bh1542_wm58_0_c20, bh1542_wm58_0_c21 :  std_logic;
signal bh1542_wm57_0_c20, bh1542_wm57_0_c21 :  std_logic;
signal bh1542_wm56_0_c20, bh1542_wm56_0_c21 :  std_logic;
signal bh1542_wm55_0_c20, bh1542_wm55_0_c21 :  std_logic;
signal bh1542_wm54_0_c20, bh1542_wm54_0_c21 :  std_logic;
signal bh1542_wm53_0_c20, bh1542_wm53_0_c21 :  std_logic;
signal bh1542_wm52_0_c20, bh1542_wm52_0_c21 :  std_logic;
signal bh1542_wm51_0_c20, bh1542_wm51_0_c21 :  std_logic;
signal bh1542_wm50_0_c20, bh1542_wm50_0_c21 :  std_logic;
signal bh1542_wm49_0_c20, bh1542_wm49_0_c21 :  std_logic;
signal bh1542_wm48_0_c20 :  std_logic;
signal bh1542_wm47_0_c20 :  std_logic;
signal bh1542_wm46_0_c20 :  std_logic;
signal bh1542_wm45_0_c20 :  std_logic;
signal bh1542_wm44_0_c20 :  std_logic;
signal bh1542_wm43_0_c20 :  std_logic;
signal bh1542_wm42_0_c20 :  std_logic;
signal bh1542_wm41_0_c20 :  std_logic;
signal bh1542_wm40_0_c20 :  std_logic;
signal bh1542_wm39_0_c20 :  std_logic;
signal bh1542_wm38_0_c20 :  std_logic;
signal bh1542_wm37_0_c20 :  std_logic;
signal bh1542_wm36_0_c20 :  std_logic;
signal bh1542_wm35_0_c20 :  std_logic;
signal bh1542_wm34_0_c20 :  std_logic;
signal bh1542_wm33_0_c20 :  std_logic;
signal bh1542_wm32_0_c20 :  std_logic;
signal bh1542_wm31_0_c20 :  std_logic;
signal bh1542_wm30_0_c20 :  std_logic;
signal bh1542_wm29_0_c20 :  std_logic;
signal bh1542_wm28_0_c20 :  std_logic;
signal bh1542_wm27_0_c20 :  std_logic;
signal bh1542_wm26_0_c20 :  std_logic;
signal bh1542_wm25_0_c20 :  std_logic;
signal tile_1_X_c19 :  std_logic_vector(1 downto 0);
signal tile_1_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_1_output_c19 :  std_logic_vector(3 downto 0);
signal tile_1_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm20_0_c19 :  std_logic;
signal bh1542_wm19_0_c19 :  std_logic;
signal bh1542_wm18_0_c19 :  std_logic;
signal bh1542_wm17_0_c19 :  std_logic;
signal tile_2_X_c19 :  std_logic_vector(2 downto 0);
signal tile_2_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_2_output_c19 :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm23_0_c19 :  std_logic;
signal bh1542_wm22_0_c19 :  std_logic;
signal bh1542_wm21_0_c19 :  std_logic;
signal bh1542_wm20_1_c19 :  std_logic;
signal bh1542_wm19_1_c19 :  std_logic;
signal tile_3_X_c19 :  std_logic_vector(2 downto 0);
signal tile_3_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_3_output_c19 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm26_1_c19, bh1542_wm26_1_c20 :  std_logic;
signal bh1542_wm25_1_c19 :  std_logic;
signal bh1542_wm24_0_c19 :  std_logic;
signal bh1542_wm23_1_c19 :  std_logic;
signal bh1542_wm22_1_c19 :  std_logic;
signal tile_4_X_c19 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_4_output_c19 :  std_logic_vector(3 downto 0);
signal tile_4_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm22_2_c19 :  std_logic;
signal bh1542_wm21_1_c19 :  std_logic;
signal bh1542_wm20_2_c19 :  std_logic;
signal bh1542_wm19_2_c19 :  std_logic;
signal tile_5_X_c19 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_5_output_c19 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm25_2_c19 :  std_logic;
signal bh1542_wm24_1_c19 :  std_logic;
signal bh1542_wm23_2_c19 :  std_logic;
signal bh1542_wm22_3_c19 :  std_logic;
signal bh1542_wm21_2_c19 :  std_logic;
signal tile_6_X_c19 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_6_output_c19 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm28_1_c19, bh1542_wm28_1_c20 :  std_logic;
signal bh1542_wm27_1_c19 :  std_logic;
signal bh1542_wm26_2_c19, bh1542_wm26_2_c20 :  std_logic;
signal bh1542_wm25_3_c19 :  std_logic;
signal bh1542_wm24_2_c19 :  std_logic;
signal tile_7_X_c19 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_7_output_c19 :  std_logic_vector(3 downto 0);
signal tile_7_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm24_3_c19 :  std_logic;
signal bh1542_wm23_3_c19 :  std_logic;
signal bh1542_wm22_4_c19 :  std_logic;
signal bh1542_wm21_3_c19 :  std_logic;
signal tile_8_X_c19 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_8_output_c19 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm27_2_c19 :  std_logic;
signal bh1542_wm26_3_c19, bh1542_wm26_3_c20 :  std_logic;
signal bh1542_wm25_4_c19 :  std_logic;
signal bh1542_wm24_4_c19 :  std_logic;
signal bh1542_wm23_4_c19 :  std_logic;
signal tile_9_X_c19 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_9_output_c19 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm30_1_c19, bh1542_wm30_1_c20 :  std_logic;
signal bh1542_wm29_1_c19, bh1542_wm29_1_c20 :  std_logic;
signal bh1542_wm28_2_c19, bh1542_wm28_2_c20 :  std_logic;
signal bh1542_wm27_3_c19 :  std_logic;
signal bh1542_wm26_4_c19, bh1542_wm26_4_c20 :  std_logic;
signal tile_10_X_c19 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_10_output_c19 :  std_logic_vector(3 downto 0);
signal tile_10_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm26_5_c19, bh1542_wm26_5_c20 :  std_logic;
signal bh1542_wm25_5_c19 :  std_logic;
signal bh1542_wm24_5_c19 :  std_logic;
signal bh1542_wm23_5_c19 :  std_logic;
signal tile_11_X_c19 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_11_output_c19 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm29_2_c19, bh1542_wm29_2_c20 :  std_logic;
signal bh1542_wm28_3_c19, bh1542_wm28_3_c20 :  std_logic;
signal bh1542_wm27_4_c19 :  std_logic;
signal bh1542_wm26_6_c19 :  std_logic;
signal bh1542_wm25_6_c19 :  std_logic;
signal tile_12_X_c19 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_12_output_c19 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm32_1_c19, bh1542_wm32_1_c20 :  std_logic;
signal bh1542_wm31_1_c19 :  std_logic;
signal bh1542_wm30_2_c19, bh1542_wm30_2_c20 :  std_logic;
signal bh1542_wm29_3_c19, bh1542_wm29_3_c20 :  std_logic;
signal bh1542_wm28_4_c19, bh1542_wm28_4_c20 :  std_logic;
signal tile_13_X_c19 :  std_logic_vector(1 downto 0);
signal tile_13_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_13_output_c19 :  std_logic_vector(3 downto 0);
signal tile_13_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm28_5_c19, bh1542_wm28_5_c20 :  std_logic;
signal bh1542_wm27_5_c19 :  std_logic;
signal bh1542_wm26_7_c19 :  std_logic;
signal bh1542_wm25_7_c19 :  std_logic;
signal tile_14_X_c19 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_14_output_c19 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm31_2_c19 :  std_logic;
signal bh1542_wm30_3_c19, bh1542_wm30_3_c20 :  std_logic;
signal bh1542_wm29_4_c19, bh1542_wm29_4_c20 :  std_logic;
signal bh1542_wm28_6_c19 :  std_logic;
signal bh1542_wm27_6_c19 :  std_logic;
signal tile_15_X_c19 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_15_output_c19 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm34_1_c19, bh1542_wm34_1_c20 :  std_logic;
signal bh1542_wm33_1_c19, bh1542_wm33_1_c20 :  std_logic;
signal bh1542_wm32_2_c19, bh1542_wm32_2_c20 :  std_logic;
signal bh1542_wm31_3_c19 :  std_logic;
signal bh1542_wm30_4_c19, bh1542_wm30_4_c20 :  std_logic;
signal tile_16_X_c19 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_16_output_c19 :  std_logic_vector(3 downto 0);
signal tile_16_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm30_5_c19, bh1542_wm30_5_c20 :  std_logic;
signal bh1542_wm29_5_c19, bh1542_wm29_5_c20 :  std_logic;
signal bh1542_wm28_7_c19 :  std_logic;
signal bh1542_wm27_7_c19 :  std_logic;
signal tile_17_X_c19 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_17_output_c19 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm33_2_c19, bh1542_wm33_2_c20 :  std_logic;
signal bh1542_wm32_3_c19, bh1542_wm32_3_c20 :  std_logic;
signal bh1542_wm31_4_c19 :  std_logic;
signal bh1542_wm30_6_c19 :  std_logic;
signal bh1542_wm29_6_c19 :  std_logic;
signal tile_18_X_c19 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_18_output_c19 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm36_1_c19, bh1542_wm36_1_c20 :  std_logic;
signal bh1542_wm35_1_c19 :  std_logic;
signal bh1542_wm34_2_c19, bh1542_wm34_2_c20 :  std_logic;
signal bh1542_wm33_3_c19, bh1542_wm33_3_c20 :  std_logic;
signal bh1542_wm32_4_c19, bh1542_wm32_4_c20 :  std_logic;
signal tile_19_X_c19 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_19_output_c19 :  std_logic_vector(3 downto 0);
signal tile_19_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm32_5_c19, bh1542_wm32_5_c20 :  std_logic;
signal bh1542_wm31_5_c19 :  std_logic;
signal bh1542_wm30_7_c19 :  std_logic;
signal bh1542_wm29_7_c19 :  std_logic;
signal tile_20_X_c19 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_20_output_c19 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm35_2_c19 :  std_logic;
signal bh1542_wm34_3_c19, bh1542_wm34_3_c20 :  std_logic;
signal bh1542_wm33_4_c19, bh1542_wm33_4_c20 :  std_logic;
signal bh1542_wm32_6_c19 :  std_logic;
signal bh1542_wm31_6_c19 :  std_logic;
signal tile_21_X_c19 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_21_output_c19 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm38_1_c19 :  std_logic;
signal bh1542_wm37_1_c19, bh1542_wm37_1_c20 :  std_logic;
signal bh1542_wm36_2_c19, bh1542_wm36_2_c20 :  std_logic;
signal bh1542_wm35_3_c19 :  std_logic;
signal bh1542_wm34_4_c19, bh1542_wm34_4_c20 :  std_logic;
signal tile_22_X_c19 :  std_logic_vector(1 downto 0);
signal tile_22_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_22_output_c19 :  std_logic_vector(3 downto 0);
signal tile_22_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm34_5_c19, bh1542_wm34_5_c20 :  std_logic;
signal bh1542_wm33_5_c19, bh1542_wm33_5_c20 :  std_logic;
signal bh1542_wm32_7_c19 :  std_logic;
signal bh1542_wm31_7_c19 :  std_logic;
signal tile_23_X_c19 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_23_output_c19 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm37_2_c19, bh1542_wm37_2_c20 :  std_logic;
signal bh1542_wm36_3_c19, bh1542_wm36_3_c20 :  std_logic;
signal bh1542_wm35_4_c19 :  std_logic;
signal bh1542_wm34_6_c19 :  std_logic;
signal bh1542_wm33_6_c19 :  std_logic;
signal tile_24_X_c19 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_24_output_c19 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm40_1_c19, bh1542_wm40_1_c20 :  std_logic;
signal bh1542_wm39_1_c19 :  std_logic;
signal bh1542_wm38_2_c19 :  std_logic;
signal bh1542_wm37_3_c19, bh1542_wm37_3_c20 :  std_logic;
signal bh1542_wm36_4_c19, bh1542_wm36_4_c20 :  std_logic;
signal tile_25_X_c19 :  std_logic_vector(1 downto 0);
signal tile_25_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_25_output_c19 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm36_5_c19, bh1542_wm36_5_c20 :  std_logic;
signal bh1542_wm35_5_c19 :  std_logic;
signal bh1542_wm34_7_c19 :  std_logic;
signal bh1542_wm33_7_c19 :  std_logic;
signal tile_26_X_c19 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_26_output_c19 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm39_2_c19 :  std_logic;
signal bh1542_wm38_3_c19 :  std_logic;
signal bh1542_wm37_4_c19, bh1542_wm37_4_c20 :  std_logic;
signal bh1542_wm36_6_c19 :  std_logic;
signal bh1542_wm35_6_c19 :  std_logic;
signal tile_27_X_c19 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_27_output_c19 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm42_1_c19 :  std_logic;
signal bh1542_wm41_1_c19, bh1542_wm41_1_c20 :  std_logic;
signal bh1542_wm40_2_c19, bh1542_wm40_2_c20 :  std_logic;
signal bh1542_wm39_3_c19 :  std_logic;
signal bh1542_wm38_4_c19 :  std_logic;
signal tile_28_X_c19 :  std_logic_vector(1 downto 0);
signal tile_28_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_28_output_c19 :  std_logic_vector(3 downto 0);
signal tile_28_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm38_5_c19 :  std_logic;
signal bh1542_wm37_5_c19, bh1542_wm37_5_c20 :  std_logic;
signal bh1542_wm36_7_c19 :  std_logic;
signal bh1542_wm35_7_c19 :  std_logic;
signal tile_29_X_c19 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_29_output_c19 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm41_2_c19, bh1542_wm41_2_c20 :  std_logic;
signal bh1542_wm40_3_c19, bh1542_wm40_3_c20 :  std_logic;
signal bh1542_wm39_4_c19 :  std_logic;
signal bh1542_wm38_6_c19 :  std_logic;
signal bh1542_wm37_6_c19 :  std_logic;
signal tile_30_X_c19 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_30_output_c19 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm44_1_c19 :  std_logic;
signal bh1542_wm43_1_c19 :  std_logic;
signal bh1542_wm42_2_c19 :  std_logic;
signal bh1542_wm41_3_c19, bh1542_wm41_3_c20 :  std_logic;
signal bh1542_wm40_4_c19, bh1542_wm40_4_c20 :  std_logic;
signal tile_31_X_c19 :  std_logic_vector(1 downto 0);
signal tile_31_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_31_output_c19 :  std_logic_vector(3 downto 0);
signal tile_31_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm40_5_c19, bh1542_wm40_5_c20 :  std_logic;
signal bh1542_wm39_5_c19 :  std_logic;
signal bh1542_wm38_7_c19 :  std_logic;
signal bh1542_wm37_7_c19 :  std_logic;
signal tile_32_X_c19 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_32_output_c19 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm43_2_c19 :  std_logic;
signal bh1542_wm42_3_c19 :  std_logic;
signal bh1542_wm41_4_c19, bh1542_wm41_4_c20 :  std_logic;
signal bh1542_wm40_6_c19 :  std_logic;
signal bh1542_wm39_6_c19 :  std_logic;
signal tile_33_X_c19 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_33_output_c19 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm46_1_c19, bh1542_wm46_1_c20 :  std_logic;
signal bh1542_wm45_1_c19, bh1542_wm45_1_c20 :  std_logic;
signal bh1542_wm44_2_c19 :  std_logic;
signal bh1542_wm43_3_c19 :  std_logic;
signal bh1542_wm42_4_c19 :  std_logic;
signal tile_34_X_c19 :  std_logic_vector(1 downto 0);
signal tile_34_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_34_output_c19 :  std_logic_vector(3 downto 0);
signal tile_34_filtered_output_c19 :  signed(3-0 downto 0);
signal bh1542_wm42_5_c19 :  std_logic;
signal bh1542_wm41_5_c19, bh1542_wm41_5_c20 :  std_logic;
signal bh1542_wm40_7_c19 :  std_logic;
signal bh1542_wm39_7_c19 :  std_logic;
signal tile_35_X_c19 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_35_output_c19 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm45_2_c19, bh1542_wm45_2_c20 :  std_logic;
signal bh1542_wm44_3_c19 :  std_logic;
signal bh1542_wm43_4_c19 :  std_logic;
signal bh1542_wm42_6_c19 :  std_logic;
signal bh1542_wm41_6_c19 :  std_logic;
signal tile_36_X_c19 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c19 :  std_logic_vector(1 downto 0);
signal tile_36_output_c19 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c19 :  unsigned(4-0 downto 0);
signal bh1542_wm48_1_c19, bh1542_wm48_1_c20 :  std_logic;
signal bh1542_wm47_1_c19, bh1542_wm47_1_c20 :  std_logic;
signal bh1542_wm46_2_c19, bh1542_wm46_2_c20 :  std_logic;
signal bh1542_wm45_3_c19, bh1542_wm45_3_c20 :  std_logic;
signal bh1542_wm44_4_c19 :  std_logic;
signal tile_37_X_c19 :  std_logic_vector(0 downto 0);
signal tile_37_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_37_output_c19 :  std_logic_vector(0 downto 0);
signal tile_37_filtered_output_c19 :  signed(0-0 downto 0);
signal bh1542_wm25_8_c19 :  std_logic;
signal tile_38_X_c19 :  std_logic_vector(3 downto 0);
signal tile_38_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_38_output_c19 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c19 :  signed(4-0 downto 0);
signal bh1542_wm29_8_c19 :  std_logic;
signal bh1542_wm28_8_c19 :  std_logic;
signal bh1542_wm27_8_c19 :  std_logic;
signal bh1542_wm26_8_c19 :  std_logic;
signal bh1542_wm25_9_c19 :  std_logic;
signal tile_39_X_c19 :  std_logic_vector(3 downto 0);
signal tile_39_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_39_output_c19 :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output_c19 :  signed(4-0 downto 0);
signal bh1542_wm33_8_c19 :  std_logic;
signal bh1542_wm32_8_c19 :  std_logic;
signal bh1542_wm31_8_c19 :  std_logic;
signal bh1542_wm30_8_c19 :  std_logic;
signal bh1542_wm29_9_c19 :  std_logic;
signal tile_40_X_c19 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_40_output_c19 :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output_c19 :  signed(4-0 downto 0);
signal bh1542_wm37_8_c19 :  std_logic;
signal bh1542_wm36_8_c19 :  std_logic;
signal bh1542_wm35_8_c19 :  std_logic;
signal bh1542_wm34_8_c19 :  std_logic;
signal bh1542_wm33_9_c19 :  std_logic;
signal tile_41_X_c19 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_41_output_c19 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c19 :  signed(4-0 downto 0);
signal bh1542_wm41_7_c19 :  std_logic;
signal bh1542_wm40_8_c19 :  std_logic;
signal bh1542_wm39_8_c19 :  std_logic;
signal bh1542_wm38_8_c19 :  std_logic;
signal bh1542_wm37_9_c19 :  std_logic;
signal tile_42_X_c19 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_42_output_c19 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c19 :  signed(4-0 downto 0);
signal bh1542_wm20_3_c19 :  std_logic;
signal bh1542_wm19_3_c19 :  std_logic;
signal bh1542_wm18_1_c19 :  std_logic;
signal bh1542_wm17_1_c19 :  std_logic;
signal bh1542_wm16_0_c19 :  std_logic;
signal tile_43_X_c19 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c19 :  std_logic_vector(0 downto 0);
signal tile_43_output_c19 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c19 :  signed(4-0 downto 0);
signal bh1542_wm24_6_c19 :  std_logic;
signal bh1542_wm23_6_c19 :  std_logic;
signal bh1542_wm22_5_c19 :  std_logic;
signal bh1542_wm21_4_c19 :  std_logic;
signal bh1542_wm20_4_c19 :  std_logic;
signal bh1542_wm41_8_c19 :  std_logic;
signal bh1542_wm40_9_c19 :  std_logic;
signal bh1542_wm39_9_c19 :  std_logic;
signal bh1542_wm38_9_c19 :  std_logic;
signal bh1542_wm37_10_c19 :  std_logic;
signal bh1542_wm36_9_c19 :  std_logic;
signal bh1542_wm35_9_c19 :  std_logic;
signal bh1542_wm34_9_c19 :  std_logic;
signal bh1542_wm33_10_c19 :  std_logic;
signal bh1542_wm32_9_c19 :  std_logic;
signal bh1542_wm31_9_c19 :  std_logic;
signal bh1542_wm30_9_c19 :  std_logic;
signal bh1542_wm29_10_c19 :  std_logic;
signal bh1542_wm28_9_c19 :  std_logic;
signal bh1542_wm27_9_c19 :  std_logic;
signal bh1542_wm26_9_c19 :  std_logic;
signal bh1542_wm25_10_c19 :  std_logic;
signal bh1542_wm24_7_c19, bh1542_wm24_7_c20 :  std_logic;
signal bh1542_wm23_7_c19 :  std_logic;
signal bh1542_wm22_6_c19 :  std_logic;
signal bh1542_wm21_5_c19 :  std_logic;
signal bh1542_wm20_5_c19 :  std_logic;
signal bh1542_wm19_4_c19 :  std_logic;
signal bh1542_wm18_2_c19 :  std_logic;
signal bh1542_wm17_2_c19 :  std_logic;
signal bh1542_wm16_1_c19 :  std_logic;
signal bh1542_wm15_0_c19 :  std_logic;
signal bh1542_wm14_0_c19 :  std_logic;
signal bh1542_wm13_0_c19 :  std_logic;
signal bh1542_wm12_0_c19 :  std_logic;
signal bh1542_wm11_0_c19 :  std_logic;
signal bh1542_wm10_0_c19 :  std_logic;
signal bh1542_wm9_0_c19 :  std_logic;
signal bh1542_wm42_7_c0, bh1542_wm42_7_c1, bh1542_wm42_7_c2, bh1542_wm42_7_c3, bh1542_wm42_7_c4, bh1542_wm42_7_c5, bh1542_wm42_7_c6, bh1542_wm42_7_c7, bh1542_wm42_7_c8, bh1542_wm42_7_c9, bh1542_wm42_7_c10, bh1542_wm42_7_c11, bh1542_wm42_7_c12, bh1542_wm42_7_c13, bh1542_wm42_7_c14, bh1542_wm42_7_c15, bh1542_wm42_7_c16, bh1542_wm42_7_c17, bh1542_wm42_7_c18, bh1542_wm42_7_c19, bh1542_wm42_7_c20 :  std_logic;
signal bh1542_wm39_10_c0, bh1542_wm39_10_c1, bh1542_wm39_10_c2, bh1542_wm39_10_c3, bh1542_wm39_10_c4, bh1542_wm39_10_c5, bh1542_wm39_10_c6, bh1542_wm39_10_c7, bh1542_wm39_10_c8, bh1542_wm39_10_c9, bh1542_wm39_10_c10, bh1542_wm39_10_c11, bh1542_wm39_10_c12, bh1542_wm39_10_c13, bh1542_wm39_10_c14, bh1542_wm39_10_c15, bh1542_wm39_10_c16, bh1542_wm39_10_c17, bh1542_wm39_10_c18, bh1542_wm39_10_c19 :  std_logic;
signal bh1542_wm38_10_c0, bh1542_wm38_10_c1, bh1542_wm38_10_c2, bh1542_wm38_10_c3, bh1542_wm38_10_c4, bh1542_wm38_10_c5, bh1542_wm38_10_c6, bh1542_wm38_10_c7, bh1542_wm38_10_c8, bh1542_wm38_10_c9, bh1542_wm38_10_c10, bh1542_wm38_10_c11, bh1542_wm38_10_c12, bh1542_wm38_10_c13, bh1542_wm38_10_c14, bh1542_wm38_10_c15, bh1542_wm38_10_c16, bh1542_wm38_10_c17, bh1542_wm38_10_c18, bh1542_wm38_10_c19, bh1542_wm38_10_c20 :  std_logic;
signal bh1542_wm37_11_c0, bh1542_wm37_11_c1, bh1542_wm37_11_c2, bh1542_wm37_11_c3, bh1542_wm37_11_c4, bh1542_wm37_11_c5, bh1542_wm37_11_c6, bh1542_wm37_11_c7, bh1542_wm37_11_c8, bh1542_wm37_11_c9, bh1542_wm37_11_c10, bh1542_wm37_11_c11, bh1542_wm37_11_c12, bh1542_wm37_11_c13, bh1542_wm37_11_c14, bh1542_wm37_11_c15, bh1542_wm37_11_c16, bh1542_wm37_11_c17, bh1542_wm37_11_c18, bh1542_wm37_11_c19 :  std_logic;
signal bh1542_wm34_10_c0, bh1542_wm34_10_c1, bh1542_wm34_10_c2, bh1542_wm34_10_c3, bh1542_wm34_10_c4, bh1542_wm34_10_c5, bh1542_wm34_10_c6, bh1542_wm34_10_c7, bh1542_wm34_10_c8, bh1542_wm34_10_c9, bh1542_wm34_10_c10, bh1542_wm34_10_c11, bh1542_wm34_10_c12, bh1542_wm34_10_c13, bh1542_wm34_10_c14, bh1542_wm34_10_c15, bh1542_wm34_10_c16, bh1542_wm34_10_c17, bh1542_wm34_10_c18, bh1542_wm34_10_c19 :  std_logic;
signal bh1542_wm33_11_c0, bh1542_wm33_11_c1, bh1542_wm33_11_c2, bh1542_wm33_11_c3, bh1542_wm33_11_c4, bh1542_wm33_11_c5, bh1542_wm33_11_c6, bh1542_wm33_11_c7, bh1542_wm33_11_c8, bh1542_wm33_11_c9, bh1542_wm33_11_c10, bh1542_wm33_11_c11, bh1542_wm33_11_c12, bh1542_wm33_11_c13, bh1542_wm33_11_c14, bh1542_wm33_11_c15, bh1542_wm33_11_c16, bh1542_wm33_11_c17, bh1542_wm33_11_c18, bh1542_wm33_11_c19 :  std_logic;
signal bh1542_wm30_10_c0, bh1542_wm30_10_c1, bh1542_wm30_10_c2, bh1542_wm30_10_c3, bh1542_wm30_10_c4, bh1542_wm30_10_c5, bh1542_wm30_10_c6, bh1542_wm30_10_c7, bh1542_wm30_10_c8, bh1542_wm30_10_c9, bh1542_wm30_10_c10, bh1542_wm30_10_c11, bh1542_wm30_10_c12, bh1542_wm30_10_c13, bh1542_wm30_10_c14, bh1542_wm30_10_c15, bh1542_wm30_10_c16, bh1542_wm30_10_c17, bh1542_wm30_10_c18, bh1542_wm30_10_c19 :  std_logic;
signal bh1542_wm29_11_c0, bh1542_wm29_11_c1, bh1542_wm29_11_c2, bh1542_wm29_11_c3, bh1542_wm29_11_c4, bh1542_wm29_11_c5, bh1542_wm29_11_c6, bh1542_wm29_11_c7, bh1542_wm29_11_c8, bh1542_wm29_11_c9, bh1542_wm29_11_c10, bh1542_wm29_11_c11, bh1542_wm29_11_c12, bh1542_wm29_11_c13, bh1542_wm29_11_c14, bh1542_wm29_11_c15, bh1542_wm29_11_c16, bh1542_wm29_11_c17, bh1542_wm29_11_c18, bh1542_wm29_11_c19 :  std_logic;
signal bh1542_wm26_10_c0, bh1542_wm26_10_c1, bh1542_wm26_10_c2, bh1542_wm26_10_c3, bh1542_wm26_10_c4, bh1542_wm26_10_c5, bh1542_wm26_10_c6, bh1542_wm26_10_c7, bh1542_wm26_10_c8, bh1542_wm26_10_c9, bh1542_wm26_10_c10, bh1542_wm26_10_c11, bh1542_wm26_10_c12, bh1542_wm26_10_c13, bh1542_wm26_10_c14, bh1542_wm26_10_c15, bh1542_wm26_10_c16, bh1542_wm26_10_c17, bh1542_wm26_10_c18, bh1542_wm26_10_c19, bh1542_wm26_10_c20 :  std_logic;
signal bh1542_wm22_7_c0, bh1542_wm22_7_c1, bh1542_wm22_7_c2, bh1542_wm22_7_c3, bh1542_wm22_7_c4, bh1542_wm22_7_c5, bh1542_wm22_7_c6, bh1542_wm22_7_c7, bh1542_wm22_7_c8, bh1542_wm22_7_c9, bh1542_wm22_7_c10, bh1542_wm22_7_c11, bh1542_wm22_7_c12, bh1542_wm22_7_c13, bh1542_wm22_7_c14, bh1542_wm22_7_c15, bh1542_wm22_7_c16, bh1542_wm22_7_c17, bh1542_wm22_7_c18, bh1542_wm22_7_c19 :  std_logic;
signal bh1542_wm18_3_c0, bh1542_wm18_3_c1, bh1542_wm18_3_c2, bh1542_wm18_3_c3, bh1542_wm18_3_c4, bh1542_wm18_3_c5, bh1542_wm18_3_c6, bh1542_wm18_3_c7, bh1542_wm18_3_c8, bh1542_wm18_3_c9, bh1542_wm18_3_c10, bh1542_wm18_3_c11, bh1542_wm18_3_c12, bh1542_wm18_3_c13, bh1542_wm18_3_c14, bh1542_wm18_3_c15, bh1542_wm18_3_c16, bh1542_wm18_3_c17, bh1542_wm18_3_c18, bh1542_wm18_3_c19 :  std_logic;
signal bh1542_wm15_1_c0, bh1542_wm15_1_c1, bh1542_wm15_1_c2, bh1542_wm15_1_c3, bh1542_wm15_1_c4, bh1542_wm15_1_c5, bh1542_wm15_1_c6, bh1542_wm15_1_c7, bh1542_wm15_1_c8, bh1542_wm15_1_c9, bh1542_wm15_1_c10, bh1542_wm15_1_c11, bh1542_wm15_1_c12, bh1542_wm15_1_c13, bh1542_wm15_1_c14, bh1542_wm15_1_c15, bh1542_wm15_1_c16, bh1542_wm15_1_c17, bh1542_wm15_1_c18, bh1542_wm15_1_c19 :  std_logic;
signal bh1542_wm14_1_c0, bh1542_wm14_1_c1, bh1542_wm14_1_c2, bh1542_wm14_1_c3, bh1542_wm14_1_c4, bh1542_wm14_1_c5, bh1542_wm14_1_c6, bh1542_wm14_1_c7, bh1542_wm14_1_c8, bh1542_wm14_1_c9, bh1542_wm14_1_c10, bh1542_wm14_1_c11, bh1542_wm14_1_c12, bh1542_wm14_1_c13, bh1542_wm14_1_c14, bh1542_wm14_1_c15, bh1542_wm14_1_c16, bh1542_wm14_1_c17, bh1542_wm14_1_c18, bh1542_wm14_1_c19 :  std_logic;
signal bh1542_wm13_1_c0, bh1542_wm13_1_c1, bh1542_wm13_1_c2, bh1542_wm13_1_c3, bh1542_wm13_1_c4, bh1542_wm13_1_c5, bh1542_wm13_1_c6, bh1542_wm13_1_c7, bh1542_wm13_1_c8, bh1542_wm13_1_c9, bh1542_wm13_1_c10, bh1542_wm13_1_c11, bh1542_wm13_1_c12, bh1542_wm13_1_c13, bh1542_wm13_1_c14, bh1542_wm13_1_c15, bh1542_wm13_1_c16, bh1542_wm13_1_c17, bh1542_wm13_1_c18, bh1542_wm13_1_c19 :  std_logic;
signal bh1542_wm12_1_c0, bh1542_wm12_1_c1, bh1542_wm12_1_c2, bh1542_wm12_1_c3, bh1542_wm12_1_c4, bh1542_wm12_1_c5, bh1542_wm12_1_c6, bh1542_wm12_1_c7, bh1542_wm12_1_c8, bh1542_wm12_1_c9, bh1542_wm12_1_c10, bh1542_wm12_1_c11, bh1542_wm12_1_c12, bh1542_wm12_1_c13, bh1542_wm12_1_c14, bh1542_wm12_1_c15, bh1542_wm12_1_c16, bh1542_wm12_1_c17, bh1542_wm12_1_c18, bh1542_wm12_1_c19 :  std_logic;
signal bh1542_wm11_1_c0, bh1542_wm11_1_c1, bh1542_wm11_1_c2, bh1542_wm11_1_c3, bh1542_wm11_1_c4, bh1542_wm11_1_c5, bh1542_wm11_1_c6, bh1542_wm11_1_c7, bh1542_wm11_1_c8, bh1542_wm11_1_c9, bh1542_wm11_1_c10, bh1542_wm11_1_c11, bh1542_wm11_1_c12, bh1542_wm11_1_c13, bh1542_wm11_1_c14, bh1542_wm11_1_c15, bh1542_wm11_1_c16, bh1542_wm11_1_c17, bh1542_wm11_1_c18, bh1542_wm11_1_c19 :  std_logic;
signal bh1542_wm10_1_c0, bh1542_wm10_1_c1, bh1542_wm10_1_c2, bh1542_wm10_1_c3, bh1542_wm10_1_c4, bh1542_wm10_1_c5, bh1542_wm10_1_c6, bh1542_wm10_1_c7, bh1542_wm10_1_c8, bh1542_wm10_1_c9, bh1542_wm10_1_c10, bh1542_wm10_1_c11, bh1542_wm10_1_c12, bh1542_wm10_1_c13, bh1542_wm10_1_c14, bh1542_wm10_1_c15, bh1542_wm10_1_c16, bh1542_wm10_1_c17, bh1542_wm10_1_c18, bh1542_wm10_1_c19 :  std_logic;
signal bh1542_wm9_1_c0, bh1542_wm9_1_c1, bh1542_wm9_1_c2, bh1542_wm9_1_c3, bh1542_wm9_1_c4, bh1542_wm9_1_c5, bh1542_wm9_1_c6, bh1542_wm9_1_c7, bh1542_wm9_1_c8, bh1542_wm9_1_c9, bh1542_wm9_1_c10, bh1542_wm9_1_c11, bh1542_wm9_1_c12, bh1542_wm9_1_c13, bh1542_wm9_1_c14, bh1542_wm9_1_c15, bh1542_wm9_1_c16, bh1542_wm9_1_c17, bh1542_wm9_1_c18, bh1542_wm9_1_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1760_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1760_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm48_2_c20, bh1542_wm48_2_c21 :  std_logic;
signal bh1542_wm47_2_c20, bh1542_wm47_2_c21 :  std_logic;
signal bh1542_wm46_3_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_copy1761_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1764_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm46_4_c20 :  std_logic;
signal bh1542_wm45_4_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_copy1765_c20 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1768_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1768_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm45_5_c20 :  std_logic;
signal bh1542_wm44_5_c20 :  std_logic;
signal bh1542_wm43_5_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_copy1769_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm44_6_c20 :  std_logic;
signal bh1542_wm43_6_c20 :  std_logic;
signal bh1542_wm42_8_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_copy1771_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm43_7_c20 :  std_logic;
signal bh1542_wm42_9_c20 :  std_logic;
signal bh1542_wm41_9_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_copy1773_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1776_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm42_10_c19, bh1542_wm42_10_c20 :  std_logic;
signal bh1542_wm41_10_c19, bh1542_wm41_10_c20 :  std_logic;
signal bh1542_wm40_10_c19, bh1542_wm40_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_copy1777_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1778_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm41_11_c20 :  std_logic;
signal bh1542_wm40_11_c20 :  std_logic;
signal bh1542_wm39_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_copy1779_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1780_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm41_12_c19, bh1542_wm41_12_c20 :  std_logic;
signal bh1542_wm40_12_c19, bh1542_wm40_12_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_copy1781_c19 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1782_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm40_13_c20 :  std_logic;
signal bh1542_wm39_12_c20 :  std_logic;
signal bh1542_wm38_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_copy1783_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm40_14_c20 :  std_logic;
signal bh1542_wm39_13_c20 :  std_logic;
signal bh1542_wm38_12_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_copy1785_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1786_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm39_14_c19, bh1542_wm39_14_c20 :  std_logic;
signal bh1542_wm38_13_c19, bh1542_wm38_13_c20 :  std_logic;
signal bh1542_wm37_12_c19, bh1542_wm37_12_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_copy1787_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm39_15_c20 :  std_logic;
signal bh1542_wm38_14_c20 :  std_logic;
signal bh1542_wm37_13_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_copy1789_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1790_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm38_15_c19, bh1542_wm38_15_c20 :  std_logic;
signal bh1542_wm37_14_c19, bh1542_wm37_14_c20 :  std_logic;
signal bh1542_wm36_10_c19, bh1542_wm36_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_copy1791_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1792_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm38_16_c19 :  std_logic;
signal bh1542_wm37_15_c19, bh1542_wm37_15_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_copy1793_c19 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1794_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm37_16_c20 :  std_logic;
signal bh1542_wm36_11_c20 :  std_logic;
signal bh1542_wm35_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_copy1795_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1796_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm37_17_c19, bh1542_wm37_17_c20 :  std_logic;
signal bh1542_wm36_12_c19, bh1542_wm36_12_c20 :  std_logic;
signal bh1542_wm35_11_c19, bh1542_wm35_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_copy1797_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1798_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm36_13_c20 :  std_logic;
signal bh1542_wm35_12_c20 :  std_logic;
signal bh1542_wm34_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_copy1799_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm36_14_c20 :  std_logic;
signal bh1542_wm35_13_c20 :  std_logic;
signal bh1542_wm34_12_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_copy1801_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1802_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm35_14_c19, bh1542_wm35_14_c20 :  std_logic;
signal bh1542_wm34_13_c19, bh1542_wm34_13_c20 :  std_logic;
signal bh1542_wm33_12_c19, bh1542_wm33_12_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_copy1803_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1804_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm35_15_c19, bh1542_wm35_15_c20 :  std_logic;
signal bh1542_wm34_14_c19, bh1542_wm34_14_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_copy1805_c19 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1806_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm34_15_c20 :  std_logic;
signal bh1542_wm33_13_c20 :  std_logic;
signal bh1542_wm32_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_copy1807_c20 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1810_In0_c19 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm34_16_c19, bh1542_wm34_16_c20 :  std_logic;
signal bh1542_wm33_14_c19, bh1542_wm33_14_c20 :  std_logic;
signal bh1542_wm32_11_c19, bh1542_wm32_11_c20 :  std_logic;
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_copy1811_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1812_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm33_15_c20 :  std_logic;
signal bh1542_wm32_12_c20 :  std_logic;
signal bh1542_wm31_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_copy1813_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1814_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm33_16_c19, bh1542_wm33_16_c20 :  std_logic;
signal bh1542_wm32_13_c19, bh1542_wm32_13_c20 :  std_logic;
signal bh1542_wm31_11_c19, bh1542_wm31_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_copy1815_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1816_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm32_14_c20 :  std_logic;
signal bh1542_wm31_12_c20 :  std_logic;
signal bh1542_wm30_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_copy1817_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm32_15_c20 :  std_logic;
signal bh1542_wm31_13_c20 :  std_logic;
signal bh1542_wm30_12_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_copy1819_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1820_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm31_14_c19, bh1542_wm31_14_c20 :  std_logic;
signal bh1542_wm30_13_c19, bh1542_wm30_13_c20 :  std_logic;
signal bh1542_wm29_12_c19, bh1542_wm29_12_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_copy1821_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1822_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm31_15_c19, bh1542_wm31_15_c20 :  std_logic;
signal bh1542_wm30_14_c19, bh1542_wm30_14_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_copy1823_c19 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1824_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm30_15_c20 :  std_logic;
signal bh1542_wm29_13_c20 :  std_logic;
signal bh1542_wm28_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_copy1825_c20 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1826_In0_c19 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm30_16_c19, bh1542_wm30_16_c20 :  std_logic;
signal bh1542_wm29_14_c19, bh1542_wm29_14_c20 :  std_logic;
signal bh1542_wm28_11_c19, bh1542_wm28_11_c20 :  std_logic;
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_copy1827_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1828_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm29_15_c20 :  std_logic;
signal bh1542_wm28_12_c20 :  std_logic;
signal bh1542_wm27_10_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_copy1829_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1830_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm29_16_c19, bh1542_wm29_16_c20 :  std_logic;
signal bh1542_wm28_13_c19, bh1542_wm28_13_c20 :  std_logic;
signal bh1542_wm27_11_c19, bh1542_wm27_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_copy1831_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1832_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm28_14_c20 :  std_logic;
signal bh1542_wm27_12_c20 :  std_logic;
signal bh1542_wm26_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_copy1833_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm28_15_c20 :  std_logic;
signal bh1542_wm27_13_c20 :  std_logic;
signal bh1542_wm26_12_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_copy1835_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1836_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm27_14_c19, bh1542_wm27_14_c20 :  std_logic;
signal bh1542_wm26_13_c19, bh1542_wm26_13_c20 :  std_logic;
signal bh1542_wm25_11_c19, bh1542_wm25_11_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_copy1837_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1838_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm27_15_c19, bh1542_wm27_15_c20 :  std_logic;
signal bh1542_wm26_14_c19, bh1542_wm26_14_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_copy1839_c19 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1840_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm26_15_c20 :  std_logic;
signal bh1542_wm25_12_c20 :  std_logic;
signal bh1542_wm24_8_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_copy1841_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In0_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm26_16_c20 :  std_logic;
signal bh1542_wm25_13_c20 :  std_logic;
signal bh1542_wm24_9_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_copy1843_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1844_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm25_14_c19, bh1542_wm25_14_c20 :  std_logic;
signal bh1542_wm24_10_c19, bh1542_wm24_10_c20 :  std_logic;
signal bh1542_wm23_8_c19 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_copy1845_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1846_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1846_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm25_15_c19, bh1542_wm25_15_c20 :  std_logic;
signal bh1542_wm24_11_c19, bh1542_wm24_11_c20 :  std_logic;
signal bh1542_wm23_9_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_copy1847_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1848_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm24_12_c19, bh1542_wm24_12_c20 :  std_logic;
signal bh1542_wm23_10_c19 :  std_logic;
signal bh1542_wm22_8_c19 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_copy1849_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1850_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm23_11_c19 :  std_logic;
signal bh1542_wm22_9_c19 :  std_logic;
signal bh1542_wm21_6_c19 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_copy1851_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1852_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1852_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm23_12_c19, bh1542_wm23_12_c20 :  std_logic;
signal bh1542_wm22_10_c19 :  std_logic;
signal bh1542_wm21_7_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_copy1853_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1854_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm22_11_c19 :  std_logic;
signal bh1542_wm21_8_c19 :  std_logic;
signal bh1542_wm20_6_c19 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_copy1855_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1856_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm21_9_c19 :  std_logic;
signal bh1542_wm20_7_c19 :  std_logic;
signal bh1542_wm19_5_c19 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_copy1857_c19 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1858_In0_c19 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm20_8_c19 :  std_logic;
signal bh1542_wm19_6_c19 :  std_logic;
signal bh1542_wm18_4_c19 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_copy1859_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1860_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1860_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm19_7_c19 :  std_logic;
signal bh1542_wm18_5_c19 :  std_logic;
signal bh1542_wm17_3_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_copy1861_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1862_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1862_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm18_6_c19 :  std_logic;
signal bh1542_wm17_4_c19 :  std_logic;
signal bh1542_wm16_2_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_copy1863_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1864_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1864_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm16_3_c19 :  std_logic;
signal bh1542_wm15_2_c19 :  std_logic;
signal bh1542_wm14_2_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_copy1865_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1866_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1866_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm14_3_c19 :  std_logic;
signal bh1542_wm13_2_c19 :  std_logic;
signal bh1542_wm12_2_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_copy1867_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1868_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1868_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm12_3_c19 :  std_logic;
signal bh1542_wm11_2_c19 :  std_logic;
signal bh1542_wm10_2_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_copy1869_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1870_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1870_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm10_3_c19 :  std_logic;
signal bh1542_wm9_2_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_copy1871_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1872_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1872_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm46_5_c20, bh1542_wm46_5_c21 :  std_logic;
signal bh1542_wm45_6_c20, bh1542_wm45_6_c21 :  std_logic;
signal bh1542_wm44_7_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_copy1873_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1874_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm44_8_c20 :  std_logic;
signal bh1542_wm43_8_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_copy1875_c20 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1876_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm43_9_c20 :  std_logic;
signal bh1542_wm42_11_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_copy1877_c20 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1878_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1878_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm42_12_c20 :  std_logic;
signal bh1542_wm41_13_c20 :  std_logic;
signal bh1542_wm40_15_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_copy1879_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1880_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm41_14_c20 :  std_logic;
signal bh1542_wm40_16_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_copy1881_c20 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1882_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1882_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm40_17_c20 :  std_logic;
signal bh1542_wm39_16_c20 :  std_logic;
signal bh1542_wm38_17_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_copy1883_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In1_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm39_17_c20 :  std_logic;
signal bh1542_wm38_18_c20 :  std_logic;
signal bh1542_wm37_18_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_copy1885_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1886_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm38_19_c20 :  std_logic;
signal bh1542_wm37_19_c20 :  std_logic;
signal bh1542_wm36_15_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_copy1887_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1888_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm37_20_c20 :  std_logic;
signal bh1542_wm36_16_c20 :  std_logic;
signal bh1542_wm35_16_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_copy1889_c20 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1890_In0_c20 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm36_17_c20 :  std_logic;
signal bh1542_wm35_17_c20 :  std_logic;
signal bh1542_wm34_17_c20 :  std_logic;
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_copy1891_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1892_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm35_18_c20 :  std_logic;
signal bh1542_wm34_18_c20 :  std_logic;
signal bh1542_wm33_17_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_copy1893_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1894_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm34_19_c20 :  std_logic;
signal bh1542_wm33_18_c20 :  std_logic;
signal bh1542_wm32_16_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_copy1895_c20 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1896_In0_c20 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm33_19_c20 :  std_logic;
signal bh1542_wm32_17_c20 :  std_logic;
signal bh1542_wm31_16_c20 :  std_logic;
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_copy1897_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1898_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm32_18_c20 :  std_logic;
signal bh1542_wm31_17_c20 :  std_logic;
signal bh1542_wm30_17_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_copy1899_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1900_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm31_18_c20 :  std_logic;
signal bh1542_wm30_18_c20 :  std_logic;
signal bh1542_wm29_17_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_copy1901_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1902_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm30_19_c20 :  std_logic;
signal bh1542_wm29_18_c20 :  std_logic;
signal bh1542_wm28_16_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_copy1903_c20 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1904_In0_c20 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm29_19_c20 :  std_logic;
signal bh1542_wm28_17_c20 :  std_logic;
signal bh1542_wm27_16_c20 :  std_logic;
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_copy1905_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1906_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm28_18_c20 :  std_logic;
signal bh1542_wm27_17_c20 :  std_logic;
signal bh1542_wm26_17_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_copy1907_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1908_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm27_18_c20 :  std_logic;
signal bh1542_wm26_18_c20 :  std_logic;
signal bh1542_wm25_16_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_copy1909_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1910_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm26_19_c20 :  std_logic;
signal bh1542_wm25_17_c20 :  std_logic;
signal bh1542_wm24_13_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_copy1911_c20 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1912_In0_c20 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm25_18_c20 :  std_logic;
signal bh1542_wm24_14_c20 :  std_logic;
signal bh1542_wm23_13_c20 :  std_logic;
signal Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_copy1913_c20 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1914_In0_c20 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm24_15_c20 :  std_logic;
signal bh1542_wm23_14_c20 :  std_logic;
signal bh1542_wm22_12_c20 :  std_logic;
signal Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_copy1915_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1916_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1916_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm23_15_c19, bh1542_wm23_15_c20 :  std_logic;
signal bh1542_wm22_13_c19, bh1542_wm22_13_c20 :  std_logic;
signal bh1542_wm21_10_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_copy1917_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1918_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm22_14_c19, bh1542_wm22_14_c20 :  std_logic;
signal bh1542_wm21_11_c19 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_copy1919_c19 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c0, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c1, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c2, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c3, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c4, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c5, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c6, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c7, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c8, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c9, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c10, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c11, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c12, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c13, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c14, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c15, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c16, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c17, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c18, Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm21_12_c19 :  std_logic;
signal bh1542_wm20_9_c19 :  std_logic;
signal bh1542_wm19_8_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_copy1921_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1922_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm20_10_c19 :  std_logic;
signal bh1542_wm19_9_c19 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_copy1923_c19 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c0, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c1, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c2, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c3, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c4, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c5, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c6, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c7, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c8, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c9, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c10, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c11, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c12, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c13, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c14, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c15, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c16, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c17, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c18, Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm19_10_c19 :  std_logic;
signal bh1542_wm18_7_c19 :  std_logic;
signal bh1542_wm17_5_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_copy1925_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1926_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_c19 :  std_logic_vector(1 downto 0);
signal bh1542_wm18_8_c19 :  std_logic;
signal bh1542_wm17_6_c19 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_copy1927_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1928_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1928_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm17_7_c19 :  std_logic;
signal bh1542_wm16_4_c19, bh1542_wm16_4_c20 :  std_logic;
signal bh1542_wm15_3_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_copy1929_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1930_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1930_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm14_4_c19 :  std_logic;
signal bh1542_wm13_3_c19, bh1542_wm13_3_c20 :  std_logic;
signal bh1542_wm12_4_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_copy1931_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1932_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1932_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm12_5_c19 :  std_logic;
signal bh1542_wm11_3_c19 :  std_logic;
signal bh1542_wm10_4_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_copy1933_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1934_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1934_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm10_5_c19 :  std_logic;
signal bh1542_wm9_3_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_copy1935_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1936_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1936_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm44_9_c20, bh1542_wm44_9_c21 :  std_logic;
signal bh1542_wm43_10_c20, bh1542_wm43_10_c21 :  std_logic;
signal bh1542_wm42_13_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_copy1937_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1938_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1938_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm42_14_c20 :  std_logic;
signal bh1542_wm41_15_c20 :  std_logic;
signal bh1542_wm40_18_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_copy1939_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1940_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1940_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm40_19_c20 :  std_logic;
signal bh1542_wm39_18_c20 :  std_logic;
signal bh1542_wm38_20_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_copy1941_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1942_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1942_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm38_21_c20 :  std_logic;
signal bh1542_wm37_21_c20 :  std_logic;
signal bh1542_wm36_18_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_copy1943_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1944_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1944_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm36_19_c20 :  std_logic;
signal bh1542_wm35_19_c20 :  std_logic;
signal bh1542_wm34_20_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_copy1945_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1946_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1946_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm34_21_c20 :  std_logic;
signal bh1542_wm33_20_c20 :  std_logic;
signal bh1542_wm32_19_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_copy1947_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1948_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1948_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm32_20_c20 :  std_logic;
signal bh1542_wm31_19_c20 :  std_logic;
signal bh1542_wm30_20_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_copy1949_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1950_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1950_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm30_21_c20 :  std_logic;
signal bh1542_wm29_20_c20 :  std_logic;
signal bh1542_wm28_19_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_copy1951_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1952_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1952_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm28_20_c20 :  std_logic;
signal bh1542_wm27_19_c20 :  std_logic;
signal bh1542_wm26_20_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_copy1953_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c0, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c1, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c2, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c3, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c4, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c5, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c6, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c7, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c8, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c9, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c10, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c11, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c12, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c13, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c14, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c15, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c16, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c17, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c18, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm26_21_c20 :  std_logic;
signal bh1542_wm25_19_c20 :  std_logic;
signal bh1542_wm24_16_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_copy1955_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1956_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm25_20_c20 :  std_logic;
signal bh1542_wm24_17_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_copy1957_c20 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1958_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm24_18_c20 :  std_logic;
signal bh1542_wm23_16_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_copy1959_c20 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c0, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c1, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c2, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c3, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c4, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c5, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c6, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c7, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c8, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c9, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c10, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c11, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c12, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c13, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c14, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c15, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c16, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c17, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c18, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm23_17_c20 :  std_logic;
signal bh1542_wm22_15_c20 :  std_logic;
signal bh1542_wm21_13_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_copy1961_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1962_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm22_16_c20 :  std_logic;
signal bh1542_wm21_14_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_copy1963_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1964_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1964_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm21_15_c20 :  std_logic;
signal bh1542_wm20_11_c20, bh1542_wm20_11_c21 :  std_logic;
signal bh1542_wm19_11_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_copy1965_c19, Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_copy1965_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1966_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1966_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm19_12_c20 :  std_logic;
signal bh1542_wm18_9_c20 :  std_logic;
signal bh1542_wm17_8_c20 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_copy1967_c19, Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_copy1967_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1968_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_c20 :  std_logic_vector(1 downto 0);
signal bh1542_wm17_9_c20 :  std_logic;
signal bh1542_wm16_5_c20 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_copy1969_c19, Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_copy1969_c20 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1970_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1970_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm15_4_c20, bh1542_wm15_4_c21 :  std_logic;
signal bh1542_wm14_5_c20, bh1542_wm14_5_c21 :  std_logic;
signal bh1542_wm13_4_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_copy1971_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_copy1971_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1972_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1972_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm12_6_c20 :  std_logic;
signal bh1542_wm11_4_c20, bh1542_wm11_4_c21 :  std_logic;
signal bh1542_wm10_6_c20 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_copy1973_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_copy1973_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1974_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1974_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh1542_wm10_7_c19, bh1542_wm10_7_c20 :  std_logic;
signal bh1542_wm9_4_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_copy1975_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1976_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1976_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm42_15_c21 :  std_logic;
signal bh1542_wm41_16_c21 :  std_logic;
signal bh1542_wm40_20_c21 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_copy1977_c20, Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_copy1977_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1978_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1978_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm40_21_c21 :  std_logic;
signal bh1542_wm39_19_c21 :  std_logic;
signal bh1542_wm38_22_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_copy1979_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_copy1979_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1980_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1980_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm38_23_c21 :  std_logic;
signal bh1542_wm37_22_c21 :  std_logic;
signal bh1542_wm36_20_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_copy1981_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_copy1981_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1982_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1982_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm36_21_c21 :  std_logic;
signal bh1542_wm35_20_c21 :  std_logic;
signal bh1542_wm34_22_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_copy1983_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_copy1983_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1984_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1984_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm34_23_c21 :  std_logic;
signal bh1542_wm33_21_c21 :  std_logic;
signal bh1542_wm32_21_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_copy1985_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_copy1985_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1986_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1986_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm32_22_c21 :  std_logic;
signal bh1542_wm31_20_c21 :  std_logic;
signal bh1542_wm30_22_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_copy1987_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_copy1987_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1988_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1988_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm30_23_c21 :  std_logic;
signal bh1542_wm29_21_c21 :  std_logic;
signal bh1542_wm28_21_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_copy1989_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_copy1989_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1990_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1990_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm28_22_c21 :  std_logic;
signal bh1542_wm27_20_c21 :  std_logic;
signal bh1542_wm26_22_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_copy1991_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_copy1991_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1992_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1992_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm26_23_c21 :  std_logic;
signal bh1542_wm25_21_c21 :  std_logic;
signal bh1542_wm24_19_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_copy1993_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_copy1993_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1994_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1994_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh1542_wm24_20_c21 :  std_logic;
signal bh1542_wm23_18_c21 :  std_logic;
signal bh1542_wm22_17_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_copy1995_c20, Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_copy1995_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1996_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_c21 :  std_logic_vector(1 downto 0);
signal bh1542_wm22_18_c21 :  std_logic;
signal bh1542_wm21_16_c21 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_copy1997_c20, Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_copy1997_c21 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1998_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_c21 :  std_logic_vector(1 downto 0);
signal bh1542_wm21_17_c21 :  std_logic;
signal bh1542_wm20_12_c21 :  std_logic;
signal Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_copy1999_c20, Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_copy1999_c21 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2000_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2000_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm19_13_c20, bh1542_wm19_13_c21 :  std_logic;
signal bh1542_wm18_10_c20, bh1542_wm18_10_c21 :  std_logic;
signal bh1542_wm17_10_c20, bh1542_wm17_10_c21 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_copy2001_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid2002_In0_c20 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid2002_In1_c20 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm17_11_c20, bh1542_wm17_11_c21 :  std_logic;
signal bh1542_wm16_6_c20, bh1542_wm16_6_c21 :  std_logic;
signal bh1542_wm15_5_c20, bh1542_wm15_5_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_copy2003_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2004_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2004_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm13_5_c20, bh1542_wm13_5_c21 :  std_logic;
signal bh1542_wm12_7_c20, bh1542_wm12_7_c21 :  std_logic;
signal bh1542_wm11_5_c20, bh1542_wm11_5_c21 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_copy2005_c20 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In0_c20 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In1_c19, Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In1_c20 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_c20 :  std_logic_vector(2 downto 0);
signal bh1542_wm10_8_c20, bh1542_wm10_8_c21 :  std_logic;
signal bh1542_wm9_5_c20, bh1542_wm9_5_c21 :  std_logic;
signal Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_copy2007_c20 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh1542_24_c21 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh1542_In0_c21 :  std_logic_vector(32 downto 0);
signal bitheapFinalAdd_bh1542_In1_c21 :  std_logic_vector(32 downto 0);
signal bitheapFinalAdd_bh1542_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh1542_Out_c21 :  std_logic_vector(32 downto 0);
signal bitheapResult_bh1542_c21 :  std_logic_vector(56 downto 0);
signal RR_c21 :  signed(-9+41 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               bh1542_wm26_1_c20 <= bh1542_wm26_1_c19;
               bh1542_wm28_1_c20 <= bh1542_wm28_1_c19;
               bh1542_wm26_2_c20 <= bh1542_wm26_2_c19;
               bh1542_wm26_3_c20 <= bh1542_wm26_3_c19;
               bh1542_wm30_1_c20 <= bh1542_wm30_1_c19;
               bh1542_wm29_1_c20 <= bh1542_wm29_1_c19;
               bh1542_wm28_2_c20 <= bh1542_wm28_2_c19;
               bh1542_wm26_4_c20 <= bh1542_wm26_4_c19;
               bh1542_wm26_5_c20 <= bh1542_wm26_5_c19;
               bh1542_wm29_2_c20 <= bh1542_wm29_2_c19;
               bh1542_wm28_3_c20 <= bh1542_wm28_3_c19;
               bh1542_wm32_1_c20 <= bh1542_wm32_1_c19;
               bh1542_wm30_2_c20 <= bh1542_wm30_2_c19;
               bh1542_wm29_3_c20 <= bh1542_wm29_3_c19;
               bh1542_wm28_4_c20 <= bh1542_wm28_4_c19;
               bh1542_wm28_5_c20 <= bh1542_wm28_5_c19;
               bh1542_wm30_3_c20 <= bh1542_wm30_3_c19;
               bh1542_wm29_4_c20 <= bh1542_wm29_4_c19;
               bh1542_wm34_1_c20 <= bh1542_wm34_1_c19;
               bh1542_wm33_1_c20 <= bh1542_wm33_1_c19;
               bh1542_wm32_2_c20 <= bh1542_wm32_2_c19;
               bh1542_wm30_4_c20 <= bh1542_wm30_4_c19;
               bh1542_wm30_5_c20 <= bh1542_wm30_5_c19;
               bh1542_wm29_5_c20 <= bh1542_wm29_5_c19;
               bh1542_wm33_2_c20 <= bh1542_wm33_2_c19;
               bh1542_wm32_3_c20 <= bh1542_wm32_3_c19;
               bh1542_wm36_1_c20 <= bh1542_wm36_1_c19;
               bh1542_wm34_2_c20 <= bh1542_wm34_2_c19;
               bh1542_wm33_3_c20 <= bh1542_wm33_3_c19;
               bh1542_wm32_4_c20 <= bh1542_wm32_4_c19;
               bh1542_wm32_5_c20 <= bh1542_wm32_5_c19;
               bh1542_wm34_3_c20 <= bh1542_wm34_3_c19;
               bh1542_wm33_4_c20 <= bh1542_wm33_4_c19;
               bh1542_wm37_1_c20 <= bh1542_wm37_1_c19;
               bh1542_wm36_2_c20 <= bh1542_wm36_2_c19;
               bh1542_wm34_4_c20 <= bh1542_wm34_4_c19;
               bh1542_wm34_5_c20 <= bh1542_wm34_5_c19;
               bh1542_wm33_5_c20 <= bh1542_wm33_5_c19;
               bh1542_wm37_2_c20 <= bh1542_wm37_2_c19;
               bh1542_wm36_3_c20 <= bh1542_wm36_3_c19;
               bh1542_wm40_1_c20 <= bh1542_wm40_1_c19;
               bh1542_wm37_3_c20 <= bh1542_wm37_3_c19;
               bh1542_wm36_4_c20 <= bh1542_wm36_4_c19;
               bh1542_wm36_5_c20 <= bh1542_wm36_5_c19;
               bh1542_wm37_4_c20 <= bh1542_wm37_4_c19;
               bh1542_wm41_1_c20 <= bh1542_wm41_1_c19;
               bh1542_wm40_2_c20 <= bh1542_wm40_2_c19;
               bh1542_wm37_5_c20 <= bh1542_wm37_5_c19;
               bh1542_wm41_2_c20 <= bh1542_wm41_2_c19;
               bh1542_wm40_3_c20 <= bh1542_wm40_3_c19;
               bh1542_wm41_3_c20 <= bh1542_wm41_3_c19;
               bh1542_wm40_4_c20 <= bh1542_wm40_4_c19;
               bh1542_wm40_5_c20 <= bh1542_wm40_5_c19;
               bh1542_wm41_4_c20 <= bh1542_wm41_4_c19;
               bh1542_wm46_1_c20 <= bh1542_wm46_1_c19;
               bh1542_wm45_1_c20 <= bh1542_wm45_1_c19;
               bh1542_wm41_5_c20 <= bh1542_wm41_5_c19;
               bh1542_wm45_2_c20 <= bh1542_wm45_2_c19;
               bh1542_wm48_1_c20 <= bh1542_wm48_1_c19;
               bh1542_wm47_1_c20 <= bh1542_wm47_1_c19;
               bh1542_wm46_2_c20 <= bh1542_wm46_2_c19;
               bh1542_wm45_3_c20 <= bh1542_wm45_3_c19;
               bh1542_wm24_7_c20 <= bh1542_wm24_7_c19;
               bh1542_wm42_7_c20 <= bh1542_wm42_7_c19;
               bh1542_wm38_10_c20 <= bh1542_wm38_10_c19;
               bh1542_wm26_10_c20 <= bh1542_wm26_10_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In0_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In0_c19;
               bh1542_wm42_10_c20 <= bh1542_wm42_10_c19;
               bh1542_wm41_10_c20 <= bh1542_wm41_10_c19;
               bh1542_wm40_10_c20 <= bh1542_wm40_10_c19;
               bh1542_wm41_12_c20 <= bh1542_wm41_12_c19;
               bh1542_wm40_12_c20 <= bh1542_wm40_12_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In0_c19;
               bh1542_wm39_14_c20 <= bh1542_wm39_14_c19;
               bh1542_wm38_13_c20 <= bh1542_wm38_13_c19;
               bh1542_wm37_12_c20 <= bh1542_wm37_12_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In0_c19;
               bh1542_wm38_15_c20 <= bh1542_wm38_15_c19;
               bh1542_wm37_14_c20 <= bh1542_wm37_14_c19;
               bh1542_wm36_10_c20 <= bh1542_wm36_10_c19;
               bh1542_wm37_15_c20 <= bh1542_wm37_15_c19;
               bh1542_wm37_17_c20 <= bh1542_wm37_17_c19;
               bh1542_wm36_12_c20 <= bh1542_wm36_12_c19;
               bh1542_wm35_11_c20 <= bh1542_wm35_11_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In0_c19;
               bh1542_wm35_14_c20 <= bh1542_wm35_14_c19;
               bh1542_wm34_13_c20 <= bh1542_wm34_13_c19;
               bh1542_wm33_12_c20 <= bh1542_wm33_12_c19;
               bh1542_wm35_15_c20 <= bh1542_wm35_15_c19;
               bh1542_wm34_14_c20 <= bh1542_wm34_14_c19;
               bh1542_wm34_16_c20 <= bh1542_wm34_16_c19;
               bh1542_wm33_14_c20 <= bh1542_wm33_14_c19;
               bh1542_wm32_11_c20 <= bh1542_wm32_11_c19;
               bh1542_wm33_16_c20 <= bh1542_wm33_16_c19;
               bh1542_wm32_13_c20 <= bh1542_wm32_13_c19;
               bh1542_wm31_11_c20 <= bh1542_wm31_11_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In0_c19;
               bh1542_wm31_14_c20 <= bh1542_wm31_14_c19;
               bh1542_wm30_13_c20 <= bh1542_wm30_13_c19;
               bh1542_wm29_12_c20 <= bh1542_wm29_12_c19;
               bh1542_wm31_15_c20 <= bh1542_wm31_15_c19;
               bh1542_wm30_14_c20 <= bh1542_wm30_14_c19;
               bh1542_wm30_16_c20 <= bh1542_wm30_16_c19;
               bh1542_wm29_14_c20 <= bh1542_wm29_14_c19;
               bh1542_wm28_11_c20 <= bh1542_wm28_11_c19;
               bh1542_wm29_16_c20 <= bh1542_wm29_16_c19;
               bh1542_wm28_13_c20 <= bh1542_wm28_13_c19;
               bh1542_wm27_11_c20 <= bh1542_wm27_11_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In0_c19;
               bh1542_wm27_14_c20 <= bh1542_wm27_14_c19;
               bh1542_wm26_13_c20 <= bh1542_wm26_13_c19;
               bh1542_wm25_11_c20 <= bh1542_wm25_11_c19;
               bh1542_wm27_15_c20 <= bh1542_wm27_15_c19;
               bh1542_wm26_14_c20 <= bh1542_wm26_14_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In0_c19;
               bh1542_wm25_14_c20 <= bh1542_wm25_14_c19;
               bh1542_wm24_10_c20 <= bh1542_wm24_10_c19;
               bh1542_wm25_15_c20 <= bh1542_wm25_15_c19;
               bh1542_wm24_11_c20 <= bh1542_wm24_11_c19;
               bh1542_wm24_12_c20 <= bh1542_wm24_12_c19;
               bh1542_wm23_12_c20 <= bh1542_wm23_12_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In1_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In1_c19;
               bh1542_wm23_15_c20 <= bh1542_wm23_15_c19;
               bh1542_wm22_13_c20 <= bh1542_wm22_13_c19;
               bh1542_wm22_14_c20 <= bh1542_wm22_14_c19;
               bh1542_wm16_4_c20 <= bh1542_wm16_4_c19;
               bh1542_wm13_3_c20 <= bh1542_wm13_3_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c19;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_copy1965_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_copy1965_c19;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_copy1967_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_copy1967_c19;
               Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_copy1969_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_copy1969_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_copy1971_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_copy1971_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_copy1973_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_copy1973_c19;
               bh1542_wm10_7_c20 <= bh1542_wm10_7_c19;
               Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In1_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In1_c19;
            end if;
            if ce_21 = '1' then
               bh1542_wm65_0_c21 <= bh1542_wm65_0_c20;
               bh1542_wm64_0_c21 <= bh1542_wm64_0_c20;
               bh1542_wm63_0_c21 <= bh1542_wm63_0_c20;
               bh1542_wm62_0_c21 <= bh1542_wm62_0_c20;
               bh1542_wm61_0_c21 <= bh1542_wm61_0_c20;
               bh1542_wm60_0_c21 <= bh1542_wm60_0_c20;
               bh1542_wm59_0_c21 <= bh1542_wm59_0_c20;
               bh1542_wm58_0_c21 <= bh1542_wm58_0_c20;
               bh1542_wm57_0_c21 <= bh1542_wm57_0_c20;
               bh1542_wm56_0_c21 <= bh1542_wm56_0_c20;
               bh1542_wm55_0_c21 <= bh1542_wm55_0_c20;
               bh1542_wm54_0_c21 <= bh1542_wm54_0_c20;
               bh1542_wm53_0_c21 <= bh1542_wm53_0_c20;
               bh1542_wm52_0_c21 <= bh1542_wm52_0_c20;
               bh1542_wm51_0_c21 <= bh1542_wm51_0_c20;
               bh1542_wm50_0_c21 <= bh1542_wm50_0_c20;
               bh1542_wm49_0_c21 <= bh1542_wm49_0_c20;
               bh1542_wm48_2_c21 <= bh1542_wm48_2_c20;
               bh1542_wm47_2_c21 <= bh1542_wm47_2_c20;
               bh1542_wm46_5_c21 <= bh1542_wm46_5_c20;
               bh1542_wm45_6_c21 <= bh1542_wm45_6_c20;
               bh1542_wm44_9_c21 <= bh1542_wm44_9_c20;
               bh1542_wm43_10_c21 <= bh1542_wm43_10_c20;
               bh1542_wm20_11_c21 <= bh1542_wm20_11_c20;
               bh1542_wm15_4_c21 <= bh1542_wm15_4_c20;
               bh1542_wm14_5_c21 <= bh1542_wm14_5_c20;
               bh1542_wm11_4_c21 <= bh1542_wm11_4_c20;
               Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_copy1977_c21 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_copy1977_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_copy1979_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_copy1979_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_copy1981_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_copy1981_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_copy1983_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_copy1983_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_copy1985_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_copy1985_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_copy1987_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_copy1987_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_copy1989_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_copy1989_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_copy1991_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_copy1991_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_copy1993_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_copy1993_c20;
               Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_copy1995_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_copy1995_c20;
               Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_copy1997_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_copy1997_c20;
               Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_copy1999_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_copy1999_c20;
               bh1542_wm19_13_c21 <= bh1542_wm19_13_c20;
               bh1542_wm18_10_c21 <= bh1542_wm18_10_c20;
               bh1542_wm17_10_c21 <= bh1542_wm17_10_c20;
               bh1542_wm17_11_c21 <= bh1542_wm17_11_c20;
               bh1542_wm16_6_c21 <= bh1542_wm16_6_c20;
               bh1542_wm15_5_c21 <= bh1542_wm15_5_c20;
               bh1542_wm13_5_c21 <= bh1542_wm13_5_c20;
               bh1542_wm12_7_c21 <= bh1542_wm12_7_c20;
               bh1542_wm11_5_c21 <= bh1542_wm11_5_c20;
               bh1542_wm10_8_c21 <= bh1542_wm10_8_c20;
               bh1542_wm9_5_c21 <= bh1542_wm9_5_c20;
            end if;
         end if;
      end process;
XX_c19 <= signed(X);
YY_c19 <= signed(Y);
AA_c19 <= signed(A);
   tile_0_X_c19 <= X(16 downto 0);
   tile_0_Y_c19 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid1544
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 X => tile_0_X_c19,
                 Y => tile_0_Y_c19,
                 R => tile_0_output_c20);

   tile_0_filtered_output_c20 <= unsigned(tile_0_output_c20(40 downto 0));
   bh1542_wm65_0_c20 <= tile_0_filtered_output_c20(0);
   bh1542_wm64_0_c20 <= tile_0_filtered_output_c20(1);
   bh1542_wm63_0_c20 <= tile_0_filtered_output_c20(2);
   bh1542_wm62_0_c20 <= tile_0_filtered_output_c20(3);
   bh1542_wm61_0_c20 <= tile_0_filtered_output_c20(4);
   bh1542_wm60_0_c20 <= tile_0_filtered_output_c20(5);
   bh1542_wm59_0_c20 <= tile_0_filtered_output_c20(6);
   bh1542_wm58_0_c20 <= tile_0_filtered_output_c20(7);
   bh1542_wm57_0_c20 <= tile_0_filtered_output_c20(8);
   bh1542_wm56_0_c20 <= tile_0_filtered_output_c20(9);
   bh1542_wm55_0_c20 <= tile_0_filtered_output_c20(10);
   bh1542_wm54_0_c20 <= tile_0_filtered_output_c20(11);
   bh1542_wm53_0_c20 <= tile_0_filtered_output_c20(12);
   bh1542_wm52_0_c20 <= tile_0_filtered_output_c20(13);
   bh1542_wm51_0_c20 <= tile_0_filtered_output_c20(14);
   bh1542_wm50_0_c20 <= tile_0_filtered_output_c20(15);
   bh1542_wm49_0_c20 <= tile_0_filtered_output_c20(16);
   bh1542_wm48_0_c20 <= tile_0_filtered_output_c20(17);
   bh1542_wm47_0_c20 <= tile_0_filtered_output_c20(18);
   bh1542_wm46_0_c20 <= tile_0_filtered_output_c20(19);
   bh1542_wm45_0_c20 <= tile_0_filtered_output_c20(20);
   bh1542_wm44_0_c20 <= tile_0_filtered_output_c20(21);
   bh1542_wm43_0_c20 <= tile_0_filtered_output_c20(22);
   bh1542_wm42_0_c20 <= tile_0_filtered_output_c20(23);
   bh1542_wm41_0_c20 <= tile_0_filtered_output_c20(24);
   bh1542_wm40_0_c20 <= tile_0_filtered_output_c20(25);
   bh1542_wm39_0_c20 <= tile_0_filtered_output_c20(26);
   bh1542_wm38_0_c20 <= tile_0_filtered_output_c20(27);
   bh1542_wm37_0_c20 <= tile_0_filtered_output_c20(28);
   bh1542_wm36_0_c20 <= tile_0_filtered_output_c20(29);
   bh1542_wm35_0_c20 <= tile_0_filtered_output_c20(30);
   bh1542_wm34_0_c20 <= tile_0_filtered_output_c20(31);
   bh1542_wm33_0_c20 <= tile_0_filtered_output_c20(32);
   bh1542_wm32_0_c20 <= tile_0_filtered_output_c20(33);
   bh1542_wm31_0_c20 <= tile_0_filtered_output_c20(34);
   bh1542_wm30_0_c20 <= tile_0_filtered_output_c20(35);
   bh1542_wm29_0_c20 <= tile_0_filtered_output_c20(36);
   bh1542_wm28_0_c20 <= tile_0_filtered_output_c20(37);
   bh1542_wm27_0_c20 <= tile_0_filtered_output_c20(38);
   bh1542_wm26_0_c20 <= tile_0_filtered_output_c20(39);
   bh1542_wm25_0_c20 <= tile_0_filtered_output_c20(40);
   tile_1_X_c19 <= X(24 downto 23);
   tile_1_Y_c19 <= Y(23 downto 22);
   tile_1_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1546
      port map ( clk  => clk,
                 X => tile_1_X_c19,
                 Y => tile_1_Y_c19,
                 R => tile_1_output_c19);

   tile_1_filtered_output_c19 <= signed(tile_1_output_c19(3 downto 0));
   bh1542_wm20_0_c19 <= tile_1_filtered_output_c19(0);
   bh1542_wm19_0_c19 <= tile_1_filtered_output_c19(1);
   bh1542_wm18_0_c19 <= tile_1_filtered_output_c19(2);
   bh1542_wm17_0_c19 <= not tile_1_filtered_output_c19(3);
   tile_2_X_c19 <= X(22 downto 20);
   tile_2_Y_c19 <= Y(23 downto 22);
   tile_2_mult: IntMultiplierLUT_3x2_Freq300_uid1551
      port map ( clk  => clk,
                 X => tile_2_X_c19,
                 Y => tile_2_Y_c19,
                 R => tile_2_output_c19);

   tile_2_filtered_output_c19 <= unsigned(tile_2_output_c19(4 downto 0));
   bh1542_wm23_0_c19 <= tile_2_filtered_output_c19(0);
   bh1542_wm22_0_c19 <= tile_2_filtered_output_c19(1);
   bh1542_wm21_0_c19 <= tile_2_filtered_output_c19(2);
   bh1542_wm20_1_c19 <= tile_2_filtered_output_c19(3);
   bh1542_wm19_1_c19 <= tile_2_filtered_output_c19(4);
   tile_3_X_c19 <= X(19 downto 17);
   tile_3_Y_c19 <= Y(23 downto 22);
   tile_3_mult: IntMultiplierLUT_3x2_Freq300_uid1556
      port map ( clk  => clk,
                 X => tile_3_X_c19,
                 Y => tile_3_Y_c19,
                 R => tile_3_output_c19);

   tile_3_filtered_output_c19 <= unsigned(tile_3_output_c19(4 downto 0));
   bh1542_wm26_1_c19 <= tile_3_filtered_output_c19(0);
   bh1542_wm25_1_c19 <= tile_3_filtered_output_c19(1);
   bh1542_wm24_0_c19 <= tile_3_filtered_output_c19(2);
   bh1542_wm23_1_c19 <= tile_3_filtered_output_c19(3);
   bh1542_wm22_1_c19 <= tile_3_filtered_output_c19(4);
   tile_4_X_c19 <= X(24 downto 23);
   tile_4_Y_c19 <= Y(21 downto 20);
   tile_4_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1561
      port map ( clk  => clk,
                 X => tile_4_X_c19,
                 Y => tile_4_Y_c19,
                 R => tile_4_output_c19);

   tile_4_filtered_output_c19 <= signed(tile_4_output_c19(3 downto 0));
   bh1542_wm22_2_c19 <= tile_4_filtered_output_c19(0);
   bh1542_wm21_1_c19 <= tile_4_filtered_output_c19(1);
   bh1542_wm20_2_c19 <= tile_4_filtered_output_c19(2);
   bh1542_wm19_2_c19 <= not tile_4_filtered_output_c19(3);
   tile_5_X_c19 <= X(22 downto 20);
   tile_5_Y_c19 <= Y(21 downto 20);
   tile_5_mult: IntMultiplierLUT_3x2_Freq300_uid1566
      port map ( clk  => clk,
                 X => tile_5_X_c19,
                 Y => tile_5_Y_c19,
                 R => tile_5_output_c19);

   tile_5_filtered_output_c19 <= unsigned(tile_5_output_c19(4 downto 0));
   bh1542_wm25_2_c19 <= tile_5_filtered_output_c19(0);
   bh1542_wm24_1_c19 <= tile_5_filtered_output_c19(1);
   bh1542_wm23_2_c19 <= tile_5_filtered_output_c19(2);
   bh1542_wm22_3_c19 <= tile_5_filtered_output_c19(3);
   bh1542_wm21_2_c19 <= tile_5_filtered_output_c19(4);
   tile_6_X_c19 <= X(19 downto 17);
   tile_6_Y_c19 <= Y(21 downto 20);
   tile_6_mult: IntMultiplierLUT_3x2_Freq300_uid1571
      port map ( clk  => clk,
                 X => tile_6_X_c19,
                 Y => tile_6_Y_c19,
                 R => tile_6_output_c19);

   tile_6_filtered_output_c19 <= unsigned(tile_6_output_c19(4 downto 0));
   bh1542_wm28_1_c19 <= tile_6_filtered_output_c19(0);
   bh1542_wm27_1_c19 <= tile_6_filtered_output_c19(1);
   bh1542_wm26_2_c19 <= tile_6_filtered_output_c19(2);
   bh1542_wm25_3_c19 <= tile_6_filtered_output_c19(3);
   bh1542_wm24_2_c19 <= tile_6_filtered_output_c19(4);
   tile_7_X_c19 <= X(24 downto 23);
   tile_7_Y_c19 <= Y(19 downto 18);
   tile_7_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1576
      port map ( clk  => clk,
                 X => tile_7_X_c19,
                 Y => tile_7_Y_c19,
                 R => tile_7_output_c19);

   tile_7_filtered_output_c19 <= signed(tile_7_output_c19(3 downto 0));
   bh1542_wm24_3_c19 <= tile_7_filtered_output_c19(0);
   bh1542_wm23_3_c19 <= tile_7_filtered_output_c19(1);
   bh1542_wm22_4_c19 <= tile_7_filtered_output_c19(2);
   bh1542_wm21_3_c19 <= not tile_7_filtered_output_c19(3);
   tile_8_X_c19 <= X(22 downto 20);
   tile_8_Y_c19 <= Y(19 downto 18);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid1581
      port map ( clk  => clk,
                 X => tile_8_X_c19,
                 Y => tile_8_Y_c19,
                 R => tile_8_output_c19);

   tile_8_filtered_output_c19 <= unsigned(tile_8_output_c19(4 downto 0));
   bh1542_wm27_2_c19 <= tile_8_filtered_output_c19(0);
   bh1542_wm26_3_c19 <= tile_8_filtered_output_c19(1);
   bh1542_wm25_4_c19 <= tile_8_filtered_output_c19(2);
   bh1542_wm24_4_c19 <= tile_8_filtered_output_c19(3);
   bh1542_wm23_4_c19 <= tile_8_filtered_output_c19(4);
   tile_9_X_c19 <= X(19 downto 17);
   tile_9_Y_c19 <= Y(19 downto 18);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid1586
      port map ( clk  => clk,
                 X => tile_9_X_c19,
                 Y => tile_9_Y_c19,
                 R => tile_9_output_c19);

   tile_9_filtered_output_c19 <= unsigned(tile_9_output_c19(4 downto 0));
   bh1542_wm30_1_c19 <= tile_9_filtered_output_c19(0);
   bh1542_wm29_1_c19 <= tile_9_filtered_output_c19(1);
   bh1542_wm28_2_c19 <= tile_9_filtered_output_c19(2);
   bh1542_wm27_3_c19 <= tile_9_filtered_output_c19(3);
   bh1542_wm26_4_c19 <= tile_9_filtered_output_c19(4);
   tile_10_X_c19 <= X(24 downto 23);
   tile_10_Y_c19 <= Y(17 downto 16);
   tile_10_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1591
      port map ( clk  => clk,
                 X => tile_10_X_c19,
                 Y => tile_10_Y_c19,
                 R => tile_10_output_c19);

   tile_10_filtered_output_c19 <= signed(tile_10_output_c19(3 downto 0));
   bh1542_wm26_5_c19 <= tile_10_filtered_output_c19(0);
   bh1542_wm25_5_c19 <= tile_10_filtered_output_c19(1);
   bh1542_wm24_5_c19 <= tile_10_filtered_output_c19(2);
   bh1542_wm23_5_c19 <= not tile_10_filtered_output_c19(3);
   tile_11_X_c19 <= X(22 downto 20);
   tile_11_Y_c19 <= Y(17 downto 16);
   tile_11_mult: IntMultiplierLUT_3x2_Freq300_uid1596
      port map ( clk  => clk,
                 X => tile_11_X_c19,
                 Y => tile_11_Y_c19,
                 R => tile_11_output_c19);

   tile_11_filtered_output_c19 <= unsigned(tile_11_output_c19(4 downto 0));
   bh1542_wm29_2_c19 <= tile_11_filtered_output_c19(0);
   bh1542_wm28_3_c19 <= tile_11_filtered_output_c19(1);
   bh1542_wm27_4_c19 <= tile_11_filtered_output_c19(2);
   bh1542_wm26_6_c19 <= tile_11_filtered_output_c19(3);
   bh1542_wm25_6_c19 <= tile_11_filtered_output_c19(4);
   tile_12_X_c19 <= X(19 downto 17);
   tile_12_Y_c19 <= Y(17 downto 16);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid1601
      port map ( clk  => clk,
                 X => tile_12_X_c19,
                 Y => tile_12_Y_c19,
                 R => tile_12_output_c19);

   tile_12_filtered_output_c19 <= unsigned(tile_12_output_c19(4 downto 0));
   bh1542_wm32_1_c19 <= tile_12_filtered_output_c19(0);
   bh1542_wm31_1_c19 <= tile_12_filtered_output_c19(1);
   bh1542_wm30_2_c19 <= tile_12_filtered_output_c19(2);
   bh1542_wm29_3_c19 <= tile_12_filtered_output_c19(3);
   bh1542_wm28_4_c19 <= tile_12_filtered_output_c19(4);
   tile_13_X_c19 <= X(24 downto 23);
   tile_13_Y_c19 <= Y(15 downto 14);
   tile_13_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1606
      port map ( clk  => clk,
                 X => tile_13_X_c19,
                 Y => tile_13_Y_c19,
                 R => tile_13_output_c19);

   tile_13_filtered_output_c19 <= signed(tile_13_output_c19(3 downto 0));
   bh1542_wm28_5_c19 <= tile_13_filtered_output_c19(0);
   bh1542_wm27_5_c19 <= tile_13_filtered_output_c19(1);
   bh1542_wm26_7_c19 <= tile_13_filtered_output_c19(2);
   bh1542_wm25_7_c19 <= not tile_13_filtered_output_c19(3);
   tile_14_X_c19 <= X(22 downto 20);
   tile_14_Y_c19 <= Y(15 downto 14);
   tile_14_mult: IntMultiplierLUT_3x2_Freq300_uid1611
      port map ( clk  => clk,
                 X => tile_14_X_c19,
                 Y => tile_14_Y_c19,
                 R => tile_14_output_c19);

   tile_14_filtered_output_c19 <= unsigned(tile_14_output_c19(4 downto 0));
   bh1542_wm31_2_c19 <= tile_14_filtered_output_c19(0);
   bh1542_wm30_3_c19 <= tile_14_filtered_output_c19(1);
   bh1542_wm29_4_c19 <= tile_14_filtered_output_c19(2);
   bh1542_wm28_6_c19 <= tile_14_filtered_output_c19(3);
   bh1542_wm27_6_c19 <= tile_14_filtered_output_c19(4);
   tile_15_X_c19 <= X(19 downto 17);
   tile_15_Y_c19 <= Y(15 downto 14);
   tile_15_mult: IntMultiplierLUT_3x2_Freq300_uid1616
      port map ( clk  => clk,
                 X => tile_15_X_c19,
                 Y => tile_15_Y_c19,
                 R => tile_15_output_c19);

   tile_15_filtered_output_c19 <= unsigned(tile_15_output_c19(4 downto 0));
   bh1542_wm34_1_c19 <= tile_15_filtered_output_c19(0);
   bh1542_wm33_1_c19 <= tile_15_filtered_output_c19(1);
   bh1542_wm32_2_c19 <= tile_15_filtered_output_c19(2);
   bh1542_wm31_3_c19 <= tile_15_filtered_output_c19(3);
   bh1542_wm30_4_c19 <= tile_15_filtered_output_c19(4);
   tile_16_X_c19 <= X(24 downto 23);
   tile_16_Y_c19 <= Y(13 downto 12);
   tile_16_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1621
      port map ( clk  => clk,
                 X => tile_16_X_c19,
                 Y => tile_16_Y_c19,
                 R => tile_16_output_c19);

   tile_16_filtered_output_c19 <= signed(tile_16_output_c19(3 downto 0));
   bh1542_wm30_5_c19 <= tile_16_filtered_output_c19(0);
   bh1542_wm29_5_c19 <= tile_16_filtered_output_c19(1);
   bh1542_wm28_7_c19 <= tile_16_filtered_output_c19(2);
   bh1542_wm27_7_c19 <= not tile_16_filtered_output_c19(3);
   tile_17_X_c19 <= X(22 downto 20);
   tile_17_Y_c19 <= Y(13 downto 12);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid1626
      port map ( clk  => clk,
                 X => tile_17_X_c19,
                 Y => tile_17_Y_c19,
                 R => tile_17_output_c19);

   tile_17_filtered_output_c19 <= unsigned(tile_17_output_c19(4 downto 0));
   bh1542_wm33_2_c19 <= tile_17_filtered_output_c19(0);
   bh1542_wm32_3_c19 <= tile_17_filtered_output_c19(1);
   bh1542_wm31_4_c19 <= tile_17_filtered_output_c19(2);
   bh1542_wm30_6_c19 <= tile_17_filtered_output_c19(3);
   bh1542_wm29_6_c19 <= tile_17_filtered_output_c19(4);
   tile_18_X_c19 <= X(19 downto 17);
   tile_18_Y_c19 <= Y(13 downto 12);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid1631
      port map ( clk  => clk,
                 X => tile_18_X_c19,
                 Y => tile_18_Y_c19,
                 R => tile_18_output_c19);

   tile_18_filtered_output_c19 <= unsigned(tile_18_output_c19(4 downto 0));
   bh1542_wm36_1_c19 <= tile_18_filtered_output_c19(0);
   bh1542_wm35_1_c19 <= tile_18_filtered_output_c19(1);
   bh1542_wm34_2_c19 <= tile_18_filtered_output_c19(2);
   bh1542_wm33_3_c19 <= tile_18_filtered_output_c19(3);
   bh1542_wm32_4_c19 <= tile_18_filtered_output_c19(4);
   tile_19_X_c19 <= X(24 downto 23);
   tile_19_Y_c19 <= Y(11 downto 10);
   tile_19_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1636
      port map ( clk  => clk,
                 X => tile_19_X_c19,
                 Y => tile_19_Y_c19,
                 R => tile_19_output_c19);

   tile_19_filtered_output_c19 <= signed(tile_19_output_c19(3 downto 0));
   bh1542_wm32_5_c19 <= tile_19_filtered_output_c19(0);
   bh1542_wm31_5_c19 <= tile_19_filtered_output_c19(1);
   bh1542_wm30_7_c19 <= tile_19_filtered_output_c19(2);
   bh1542_wm29_7_c19 <= not tile_19_filtered_output_c19(3);
   tile_20_X_c19 <= X(22 downto 20);
   tile_20_Y_c19 <= Y(11 downto 10);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid1641
      port map ( clk  => clk,
                 X => tile_20_X_c19,
                 Y => tile_20_Y_c19,
                 R => tile_20_output_c19);

   tile_20_filtered_output_c19 <= unsigned(tile_20_output_c19(4 downto 0));
   bh1542_wm35_2_c19 <= tile_20_filtered_output_c19(0);
   bh1542_wm34_3_c19 <= tile_20_filtered_output_c19(1);
   bh1542_wm33_4_c19 <= tile_20_filtered_output_c19(2);
   bh1542_wm32_6_c19 <= tile_20_filtered_output_c19(3);
   bh1542_wm31_6_c19 <= tile_20_filtered_output_c19(4);
   tile_21_X_c19 <= X(19 downto 17);
   tile_21_Y_c19 <= Y(11 downto 10);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid1646
      port map ( clk  => clk,
                 X => tile_21_X_c19,
                 Y => tile_21_Y_c19,
                 R => tile_21_output_c19);

   tile_21_filtered_output_c19 <= unsigned(tile_21_output_c19(4 downto 0));
   bh1542_wm38_1_c19 <= tile_21_filtered_output_c19(0);
   bh1542_wm37_1_c19 <= tile_21_filtered_output_c19(1);
   bh1542_wm36_2_c19 <= tile_21_filtered_output_c19(2);
   bh1542_wm35_3_c19 <= tile_21_filtered_output_c19(3);
   bh1542_wm34_4_c19 <= tile_21_filtered_output_c19(4);
   tile_22_X_c19 <= X(24 downto 23);
   tile_22_Y_c19 <= Y(9 downto 8);
   tile_22_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1651
      port map ( clk  => clk,
                 X => tile_22_X_c19,
                 Y => tile_22_Y_c19,
                 R => tile_22_output_c19);

   tile_22_filtered_output_c19 <= signed(tile_22_output_c19(3 downto 0));
   bh1542_wm34_5_c19 <= tile_22_filtered_output_c19(0);
   bh1542_wm33_5_c19 <= tile_22_filtered_output_c19(1);
   bh1542_wm32_7_c19 <= tile_22_filtered_output_c19(2);
   bh1542_wm31_7_c19 <= not tile_22_filtered_output_c19(3);
   tile_23_X_c19 <= X(22 downto 20);
   tile_23_Y_c19 <= Y(9 downto 8);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid1656
      port map ( clk  => clk,
                 X => tile_23_X_c19,
                 Y => tile_23_Y_c19,
                 R => tile_23_output_c19);

   tile_23_filtered_output_c19 <= unsigned(tile_23_output_c19(4 downto 0));
   bh1542_wm37_2_c19 <= tile_23_filtered_output_c19(0);
   bh1542_wm36_3_c19 <= tile_23_filtered_output_c19(1);
   bh1542_wm35_4_c19 <= tile_23_filtered_output_c19(2);
   bh1542_wm34_6_c19 <= tile_23_filtered_output_c19(3);
   bh1542_wm33_6_c19 <= tile_23_filtered_output_c19(4);
   tile_24_X_c19 <= X(19 downto 17);
   tile_24_Y_c19 <= Y(9 downto 8);
   tile_24_mult: IntMultiplierLUT_3x2_Freq300_uid1661
      port map ( clk  => clk,
                 X => tile_24_X_c19,
                 Y => tile_24_Y_c19,
                 R => tile_24_output_c19);

   tile_24_filtered_output_c19 <= unsigned(tile_24_output_c19(4 downto 0));
   bh1542_wm40_1_c19 <= tile_24_filtered_output_c19(0);
   bh1542_wm39_1_c19 <= tile_24_filtered_output_c19(1);
   bh1542_wm38_2_c19 <= tile_24_filtered_output_c19(2);
   bh1542_wm37_3_c19 <= tile_24_filtered_output_c19(3);
   bh1542_wm36_4_c19 <= tile_24_filtered_output_c19(4);
   tile_25_X_c19 <= X(24 downto 23);
   tile_25_Y_c19 <= Y(7 downto 6);
   tile_25_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1666
      port map ( clk  => clk,
                 X => tile_25_X_c19,
                 Y => tile_25_Y_c19,
                 R => tile_25_output_c19);

   tile_25_filtered_output_c19 <= signed(tile_25_output_c19(3 downto 0));
   bh1542_wm36_5_c19 <= tile_25_filtered_output_c19(0);
   bh1542_wm35_5_c19 <= tile_25_filtered_output_c19(1);
   bh1542_wm34_7_c19 <= tile_25_filtered_output_c19(2);
   bh1542_wm33_7_c19 <= not tile_25_filtered_output_c19(3);
   tile_26_X_c19 <= X(22 downto 20);
   tile_26_Y_c19 <= Y(7 downto 6);
   tile_26_mult: IntMultiplierLUT_3x2_Freq300_uid1671
      port map ( clk  => clk,
                 X => tile_26_X_c19,
                 Y => tile_26_Y_c19,
                 R => tile_26_output_c19);

   tile_26_filtered_output_c19 <= unsigned(tile_26_output_c19(4 downto 0));
   bh1542_wm39_2_c19 <= tile_26_filtered_output_c19(0);
   bh1542_wm38_3_c19 <= tile_26_filtered_output_c19(1);
   bh1542_wm37_4_c19 <= tile_26_filtered_output_c19(2);
   bh1542_wm36_6_c19 <= tile_26_filtered_output_c19(3);
   bh1542_wm35_6_c19 <= tile_26_filtered_output_c19(4);
   tile_27_X_c19 <= X(19 downto 17);
   tile_27_Y_c19 <= Y(7 downto 6);
   tile_27_mult: IntMultiplierLUT_3x2_Freq300_uid1676
      port map ( clk  => clk,
                 X => tile_27_X_c19,
                 Y => tile_27_Y_c19,
                 R => tile_27_output_c19);

   tile_27_filtered_output_c19 <= unsigned(tile_27_output_c19(4 downto 0));
   bh1542_wm42_1_c19 <= tile_27_filtered_output_c19(0);
   bh1542_wm41_1_c19 <= tile_27_filtered_output_c19(1);
   bh1542_wm40_2_c19 <= tile_27_filtered_output_c19(2);
   bh1542_wm39_3_c19 <= tile_27_filtered_output_c19(3);
   bh1542_wm38_4_c19 <= tile_27_filtered_output_c19(4);
   tile_28_X_c19 <= X(24 downto 23);
   tile_28_Y_c19 <= Y(5 downto 4);
   tile_28_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1681
      port map ( clk  => clk,
                 X => tile_28_X_c19,
                 Y => tile_28_Y_c19,
                 R => tile_28_output_c19);

   tile_28_filtered_output_c19 <= signed(tile_28_output_c19(3 downto 0));
   bh1542_wm38_5_c19 <= tile_28_filtered_output_c19(0);
   bh1542_wm37_5_c19 <= tile_28_filtered_output_c19(1);
   bh1542_wm36_7_c19 <= tile_28_filtered_output_c19(2);
   bh1542_wm35_7_c19 <= not tile_28_filtered_output_c19(3);
   tile_29_X_c19 <= X(22 downto 20);
   tile_29_Y_c19 <= Y(5 downto 4);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid1686
      port map ( clk  => clk,
                 X => tile_29_X_c19,
                 Y => tile_29_Y_c19,
                 R => tile_29_output_c19);

   tile_29_filtered_output_c19 <= unsigned(tile_29_output_c19(4 downto 0));
   bh1542_wm41_2_c19 <= tile_29_filtered_output_c19(0);
   bh1542_wm40_3_c19 <= tile_29_filtered_output_c19(1);
   bh1542_wm39_4_c19 <= tile_29_filtered_output_c19(2);
   bh1542_wm38_6_c19 <= tile_29_filtered_output_c19(3);
   bh1542_wm37_6_c19 <= tile_29_filtered_output_c19(4);
   tile_30_X_c19 <= X(19 downto 17);
   tile_30_Y_c19 <= Y(5 downto 4);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid1691
      port map ( clk  => clk,
                 X => tile_30_X_c19,
                 Y => tile_30_Y_c19,
                 R => tile_30_output_c19);

   tile_30_filtered_output_c19 <= unsigned(tile_30_output_c19(4 downto 0));
   bh1542_wm44_1_c19 <= tile_30_filtered_output_c19(0);
   bh1542_wm43_1_c19 <= tile_30_filtered_output_c19(1);
   bh1542_wm42_2_c19 <= tile_30_filtered_output_c19(2);
   bh1542_wm41_3_c19 <= tile_30_filtered_output_c19(3);
   bh1542_wm40_4_c19 <= tile_30_filtered_output_c19(4);
   tile_31_X_c19 <= X(24 downto 23);
   tile_31_Y_c19 <= Y(3 downto 2);
   tile_31_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1696
      port map ( clk  => clk,
                 X => tile_31_X_c19,
                 Y => tile_31_Y_c19,
                 R => tile_31_output_c19);

   tile_31_filtered_output_c19 <= signed(tile_31_output_c19(3 downto 0));
   bh1542_wm40_5_c19 <= tile_31_filtered_output_c19(0);
   bh1542_wm39_5_c19 <= tile_31_filtered_output_c19(1);
   bh1542_wm38_7_c19 <= tile_31_filtered_output_c19(2);
   bh1542_wm37_7_c19 <= not tile_31_filtered_output_c19(3);
   tile_32_X_c19 <= X(22 downto 20);
   tile_32_Y_c19 <= Y(3 downto 2);
   tile_32_mult: IntMultiplierLUT_3x2_Freq300_uid1701
      port map ( clk  => clk,
                 X => tile_32_X_c19,
                 Y => tile_32_Y_c19,
                 R => tile_32_output_c19);

   tile_32_filtered_output_c19 <= unsigned(tile_32_output_c19(4 downto 0));
   bh1542_wm43_2_c19 <= tile_32_filtered_output_c19(0);
   bh1542_wm42_3_c19 <= tile_32_filtered_output_c19(1);
   bh1542_wm41_4_c19 <= tile_32_filtered_output_c19(2);
   bh1542_wm40_6_c19 <= tile_32_filtered_output_c19(3);
   bh1542_wm39_6_c19 <= tile_32_filtered_output_c19(4);
   tile_33_X_c19 <= X(19 downto 17);
   tile_33_Y_c19 <= Y(3 downto 2);
   tile_33_mult: IntMultiplierLUT_3x2_Freq300_uid1706
      port map ( clk  => clk,
                 X => tile_33_X_c19,
                 Y => tile_33_Y_c19,
                 R => tile_33_output_c19);

   tile_33_filtered_output_c19 <= unsigned(tile_33_output_c19(4 downto 0));
   bh1542_wm46_1_c19 <= tile_33_filtered_output_c19(0);
   bh1542_wm45_1_c19 <= tile_33_filtered_output_c19(1);
   bh1542_wm44_2_c19 <= tile_33_filtered_output_c19(2);
   bh1542_wm43_3_c19 <= tile_33_filtered_output_c19(3);
   bh1542_wm42_4_c19 <= tile_33_filtered_output_c19(4);
   tile_34_X_c19 <= X(24 downto 23);
   tile_34_Y_c19 <= Y(1 downto 0);
   tile_34_mult: IntMultiplierLUT_2_signedx2_Freq300_uid1711
      port map ( clk  => clk,
                 X => tile_34_X_c19,
                 Y => tile_34_Y_c19,
                 R => tile_34_output_c19);

   tile_34_filtered_output_c19 <= signed(tile_34_output_c19(3 downto 0));
   bh1542_wm42_5_c19 <= tile_34_filtered_output_c19(0);
   bh1542_wm41_5_c19 <= tile_34_filtered_output_c19(1);
   bh1542_wm40_7_c19 <= tile_34_filtered_output_c19(2);
   bh1542_wm39_7_c19 <= not tile_34_filtered_output_c19(3);
   tile_35_X_c19 <= X(22 downto 20);
   tile_35_Y_c19 <= Y(1 downto 0);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid1716
      port map ( clk  => clk,
                 X => tile_35_X_c19,
                 Y => tile_35_Y_c19,
                 R => tile_35_output_c19);

   tile_35_filtered_output_c19 <= unsigned(tile_35_output_c19(4 downto 0));
   bh1542_wm45_2_c19 <= tile_35_filtered_output_c19(0);
   bh1542_wm44_3_c19 <= tile_35_filtered_output_c19(1);
   bh1542_wm43_4_c19 <= tile_35_filtered_output_c19(2);
   bh1542_wm42_6_c19 <= tile_35_filtered_output_c19(3);
   bh1542_wm41_6_c19 <= tile_35_filtered_output_c19(4);
   tile_36_X_c19 <= X(19 downto 17);
   tile_36_Y_c19 <= Y(1 downto 0);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid1721
      port map ( clk  => clk,
                 X => tile_36_X_c19,
                 Y => tile_36_Y_c19,
                 R => tile_36_output_c19);

   tile_36_filtered_output_c19 <= unsigned(tile_36_output_c19(4 downto 0));
   bh1542_wm48_1_c19 <= tile_36_filtered_output_c19(0);
   bh1542_wm47_1_c19 <= tile_36_filtered_output_c19(1);
   bh1542_wm46_2_c19 <= tile_36_filtered_output_c19(2);
   bh1542_wm45_3_c19 <= tile_36_filtered_output_c19(3);
   bh1542_wm44_4_c19 <= tile_36_filtered_output_c19(4);
   tile_37_X_c19 <= X(16 downto 16);
   tile_37_Y_c19 <= Y(24 downto 24);
   tile_37_mult: IntMultiplierLUT_1x1_signed_Freq300_uid1726
      port map ( clk  => clk,
                 X => tile_37_X_c19,
                 Y => tile_37_Y_c19,
                 R => tile_37_output_c19);

   tile_37_filtered_output_c19 <= signed(tile_37_output_c19(0 downto 0));
   bh1542_wm25_8_c19 <= not tile_37_filtered_output_c19(0);
   tile_38_X_c19 <= X(15 downto 12);
   tile_38_Y_c19 <= Y(24 downto 24);
   tile_38_mult: IntMultiplierLUT_4x1_signed_Freq300_uid1728
      port map ( clk  => clk,
                 X => tile_38_X_c19,
                 Y => tile_38_Y_c19,
                 R => tile_38_output_c19);

   tile_38_filtered_output_c19 <= signed(tile_38_output_c19(4 downto 0));
   bh1542_wm29_8_c19 <= tile_38_filtered_output_c19(0);
   bh1542_wm28_8_c19 <= tile_38_filtered_output_c19(1);
   bh1542_wm27_8_c19 <= tile_38_filtered_output_c19(2);
   bh1542_wm26_8_c19 <= tile_38_filtered_output_c19(3);
   bh1542_wm25_9_c19 <= not tile_38_filtered_output_c19(4);
   tile_39_X_c19 <= X(11 downto 8);
   tile_39_Y_c19 <= Y(24 downto 24);
   tile_39_mult: IntMultiplierLUT_4x1_signed_Freq300_uid1733
      port map ( clk  => clk,
                 X => tile_39_X_c19,
                 Y => tile_39_Y_c19,
                 R => tile_39_output_c19);

   tile_39_filtered_output_c19 <= signed(tile_39_output_c19(4 downto 0));
   bh1542_wm33_8_c19 <= tile_39_filtered_output_c19(0);
   bh1542_wm32_8_c19 <= tile_39_filtered_output_c19(1);
   bh1542_wm31_8_c19 <= tile_39_filtered_output_c19(2);
   bh1542_wm30_8_c19 <= tile_39_filtered_output_c19(3);
   bh1542_wm29_9_c19 <= not tile_39_filtered_output_c19(4);
   tile_40_X_c19 <= X(7 downto 4);
   tile_40_Y_c19 <= Y(24 downto 24);
   tile_40_mult: IntMultiplierLUT_4x1_signed_Freq300_uid1738
      port map ( clk  => clk,
                 X => tile_40_X_c19,
                 Y => tile_40_Y_c19,
                 R => tile_40_output_c19);

   tile_40_filtered_output_c19 <= signed(tile_40_output_c19(4 downto 0));
   bh1542_wm37_8_c19 <= tile_40_filtered_output_c19(0);
   bh1542_wm36_8_c19 <= tile_40_filtered_output_c19(1);
   bh1542_wm35_8_c19 <= tile_40_filtered_output_c19(2);
   bh1542_wm34_8_c19 <= tile_40_filtered_output_c19(3);
   bh1542_wm33_9_c19 <= not tile_40_filtered_output_c19(4);
   tile_41_X_c19 <= X(3 downto 0);
   tile_41_Y_c19 <= Y(24 downto 24);
   tile_41_mult: IntMultiplierLUT_4x1_signed_Freq300_uid1743
      port map ( clk  => clk,
                 X => tile_41_X_c19,
                 Y => tile_41_Y_c19,
                 R => tile_41_output_c19);

   tile_41_filtered_output_c19 <= signed(tile_41_output_c19(4 downto 0));
   bh1542_wm41_7_c19 <= tile_41_filtered_output_c19(0);
   bh1542_wm40_8_c19 <= tile_41_filtered_output_c19(1);
   bh1542_wm39_8_c19 <= tile_41_filtered_output_c19(2);
   bh1542_wm38_8_c19 <= tile_41_filtered_output_c19(3);
   bh1542_wm37_9_c19 <= not tile_41_filtered_output_c19(4);
   tile_42_X_c19 <= X(24 downto 21);
   tile_42_Y_c19 <= Y(24 downto 24);
   tile_42_mult: IntMultiplierLUT_4_signedx1_signed_Freq300_uid1748
      port map ( clk  => clk,
                 X => tile_42_X_c19,
                 Y => tile_42_Y_c19,
                 R => tile_42_output_c19);

   tile_42_filtered_output_c19 <= signed(tile_42_output_c19(4 downto 0));
   bh1542_wm20_3_c19 <= tile_42_filtered_output_c19(0);
   bh1542_wm19_3_c19 <= tile_42_filtered_output_c19(1);
   bh1542_wm18_1_c19 <= tile_42_filtered_output_c19(2);
   bh1542_wm17_1_c19 <= tile_42_filtered_output_c19(3);
   bh1542_wm16_0_c19 <= not tile_42_filtered_output_c19(4);
   tile_43_X_c19 <= X(20 downto 17);
   tile_43_Y_c19 <= Y(24 downto 24);
   tile_43_mult: IntMultiplierLUT_4x1_signed_Freq300_uid1753
      port map ( clk  => clk,
                 X => tile_43_X_c19,
                 Y => tile_43_Y_c19,
                 R => tile_43_output_c19);

   tile_43_filtered_output_c19 <= signed(tile_43_output_c19(4 downto 0));
   bh1542_wm24_6_c19 <= tile_43_filtered_output_c19(0);
   bh1542_wm23_6_c19 <= tile_43_filtered_output_c19(1);
   bh1542_wm22_5_c19 <= tile_43_filtered_output_c19(2);
   bh1542_wm21_4_c19 <= tile_43_filtered_output_c19(3);
   bh1542_wm20_4_c19 <= not tile_43_filtered_output_c19(4);
   bh1542_wm41_8_c19 <= AA_c19(0);
   bh1542_wm40_9_c19 <= AA_c19(1);
   bh1542_wm39_9_c19 <= AA_c19(2);
   bh1542_wm38_9_c19 <= AA_c19(3);
   bh1542_wm37_10_c19 <= AA_c19(4);
   bh1542_wm36_9_c19 <= AA_c19(5);
   bh1542_wm35_9_c19 <= AA_c19(6);
   bh1542_wm34_9_c19 <= AA_c19(7);
   bh1542_wm33_10_c19 <= AA_c19(8);
   bh1542_wm32_9_c19 <= AA_c19(9);
   bh1542_wm31_9_c19 <= AA_c19(10);
   bh1542_wm30_9_c19 <= AA_c19(11);
   bh1542_wm29_10_c19 <= AA_c19(12);
   bh1542_wm28_9_c19 <= AA_c19(13);
   bh1542_wm27_9_c19 <= AA_c19(14);
   bh1542_wm26_9_c19 <= AA_c19(15);
   bh1542_wm25_10_c19 <= AA_c19(16);
   bh1542_wm24_7_c19 <= AA_c19(17);
   bh1542_wm23_7_c19 <= AA_c19(18);
   bh1542_wm22_6_c19 <= AA_c19(19);
   bh1542_wm21_5_c19 <= AA_c19(20);
   bh1542_wm20_5_c19 <= AA_c19(21);
   bh1542_wm19_4_c19 <= AA_c19(22);
   bh1542_wm18_2_c19 <= AA_c19(23);
   bh1542_wm17_2_c19 <= AA_c19(24);
   bh1542_wm16_1_c19 <= AA_c19(25);
   bh1542_wm15_0_c19 <= AA_c19(26);
   bh1542_wm14_0_c19 <= AA_c19(27);
   bh1542_wm13_0_c19 <= AA_c19(28);
   bh1542_wm12_0_c19 <= AA_c19(29);
   bh1542_wm11_0_c19 <= AA_c19(30);
   bh1542_wm10_0_c19 <= AA_c19(31);
   bh1542_wm9_0_c19 <= AA_c19(32);

   -- Adding the constant bits 
   bh1542_wm42_7_c0 <= '1';
   bh1542_wm39_10_c0 <= '1';
   bh1542_wm38_10_c0 <= '1';
   bh1542_wm37_11_c0 <= '1';
   bh1542_wm34_10_c0 <= '1';
   bh1542_wm33_11_c0 <= '1';
   bh1542_wm30_10_c0 <= '1';
   bh1542_wm29_11_c0 <= '1';
   bh1542_wm26_10_c0 <= '1';
   bh1542_wm22_7_c0 <= '1';
   bh1542_wm18_3_c0 <= '1';
   bh1542_wm15_1_c0 <= '1';
   bh1542_wm14_1_c0 <= '1';
   bh1542_wm13_1_c0 <= '1';
   bh1542_wm12_1_c0 <= '1';
   bh1542_wm11_1_c0 <= '1';
   bh1542_wm10_1_c0 <= '1';
   bh1542_wm9_1_c0 <= '1';


   Compressor_23_3_Freq300_uid1759_bh1542_uid1760_In0_c20 <= "" & bh1542_wm48_0_c20 & bh1542_wm48_1_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1760_In1_c20 <= "" & bh1542_wm47_0_c20 & bh1542_wm47_1_c20;
   bh1542_wm48_2_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_c20(0);
   bh1542_wm47_2_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_c20(1);
   bh1542_wm46_3_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1760: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1760_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1760_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_copy1761_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1760_Out0_copy1761_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1764_In0_c20 <= "" & bh1542_wm46_0_c20 & bh1542_wm46_1_c20 & bh1542_wm46_2_c20;
   bh1542_wm46_4_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_c20(0);
   bh1542_wm45_4_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1764: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1764_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_copy1765_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1764_Out0_copy1765_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1768_In0_c20 <= "" & bh1542_wm45_0_c20 & bh1542_wm45_1_c20 & bh1542_wm45_2_c20 & bh1542_wm45_3_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1768_In1_c20 <= "" & bh1542_wm44_0_c20;
   bh1542_wm45_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_c20(0);
   bh1542_wm44_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_c20(1);
   bh1542_wm43_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1768: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1768_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1768_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_copy1769_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1768_Out0_copy1769_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In0_c19 <= "" & bh1542_wm44_1_c19 & bh1542_wm44_2_c19 & bh1542_wm44_3_c19 & bh1542_wm44_4_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In1_c20 <= "" & bh1542_wm43_0_c20;
   bh1542_wm44_6_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_c20(0);
   bh1542_wm43_6_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_c20(1);
   bh1542_wm42_8_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1770: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1770_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_copy1771_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1770_Out0_copy1771_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In0_c19 <= "" & bh1542_wm43_1_c19 & bh1542_wm43_2_c19 & bh1542_wm43_3_c19 & bh1542_wm43_4_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In1_c20 <= "" & bh1542_wm42_0_c20;
   bh1542_wm43_7_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_c20(0);
   bh1542_wm42_9_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_c20(1);
   bh1542_wm41_9_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1772: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1772_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_copy1773_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1772_Out0_copy1773_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1776_In0_c19 <= "" & bh1542_wm42_1_c19 & bh1542_wm42_2_c19 & bh1542_wm42_3_c19 & bh1542_wm42_4_c19 & bh1542_wm42_5_c19 & bh1542_wm42_6_c19;
   bh1542_wm42_10_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_c19(0);
   bh1542_wm41_10_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_c19(1);
   bh1542_wm40_10_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1776: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1776_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_copy1777_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1776_Out0_copy1777_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1778_In0_c20 <= "" & bh1542_wm41_0_c20 & bh1542_wm41_1_c20 & bh1542_wm41_2_c20 & bh1542_wm41_3_c20 & bh1542_wm41_4_c20 & bh1542_wm41_5_c20;
   bh1542_wm41_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_c20(0);
   bh1542_wm40_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_c20(1);
   bh1542_wm39_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1778: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1778_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_copy1779_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1778_Out0_copy1779_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1780_In0_c19 <= "" & bh1542_wm41_6_c19 & bh1542_wm41_7_c19 & bh1542_wm41_8_c19;
   bh1542_wm41_12_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_c19(0);
   bh1542_wm40_12_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1780: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1780_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_copy1781_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1780_Out0_copy1781_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1782_In0_c20 <= "" & bh1542_wm40_0_c20 & bh1542_wm40_1_c20 & bh1542_wm40_2_c20 & bh1542_wm40_3_c20 & bh1542_wm40_4_c20 & bh1542_wm40_5_c20;
   bh1542_wm40_13_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_c20(0);
   bh1542_wm39_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_c20(1);
   bh1542_wm38_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1782: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1782_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_copy1783_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1782_Out0_copy1783_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In0_c19 <= "" & bh1542_wm40_6_c19 & bh1542_wm40_7_c19 & bh1542_wm40_8_c19 & bh1542_wm40_9_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In1_c20 <= "" & bh1542_wm39_0_c20;
   bh1542_wm40_14_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_c20(0);
   bh1542_wm39_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_c20(1);
   bh1542_wm38_12_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1784: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1784_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_copy1785_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1784_Out0_copy1785_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1786_In0_c19 <= "" & bh1542_wm39_1_c19 & bh1542_wm39_2_c19 & bh1542_wm39_3_c19 & bh1542_wm39_4_c19 & bh1542_wm39_5_c19 & bh1542_wm39_6_c19;
   bh1542_wm39_14_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_c19(0);
   bh1542_wm38_13_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_c19(1);
   bh1542_wm37_12_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1786: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1786_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_copy1787_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1786_Out0_copy1787_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In0_c19 <= "" & bh1542_wm39_7_c19 & bh1542_wm39_8_c19 & bh1542_wm39_9_c19 & bh1542_wm39_10_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In1_c20 <= "" & bh1542_wm38_0_c20;
   bh1542_wm39_15_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_c20(0);
   bh1542_wm38_14_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_c20(1);
   bh1542_wm37_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1788: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1788_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_copy1789_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1788_Out0_copy1789_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1790_In0_c19 <= "" & bh1542_wm38_1_c19 & bh1542_wm38_2_c19 & bh1542_wm38_3_c19 & bh1542_wm38_4_c19 & bh1542_wm38_5_c19 & bh1542_wm38_6_c19;
   bh1542_wm38_15_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_c19(0);
   bh1542_wm37_14_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_c19(1);
   bh1542_wm36_10_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1790: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1790_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_copy1791_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1790_Out0_copy1791_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1792_In0_c19 <= "" & bh1542_wm38_7_c19 & bh1542_wm38_8_c19 & bh1542_wm38_9_c19;
   bh1542_wm38_16_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_c19(0);
   bh1542_wm37_15_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1792: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1792_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_copy1793_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1792_Out0_copy1793_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1794_In0_c20 <= "" & bh1542_wm37_0_c20 & bh1542_wm37_1_c20 & bh1542_wm37_2_c20 & bh1542_wm37_3_c20 & bh1542_wm37_4_c20 & bh1542_wm37_5_c20;
   bh1542_wm37_16_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_c20(0);
   bh1542_wm36_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_c20(1);
   bh1542_wm35_10_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1794: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1794_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_copy1795_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1794_Out0_copy1795_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1796_In0_c19 <= "" & bh1542_wm37_8_c19 & bh1542_wm37_11_c19 & bh1542_wm37_10_c19 & bh1542_wm37_9_c19 & bh1542_wm37_7_c19 & bh1542_wm37_6_c19;
   bh1542_wm37_17_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_c19(0);
   bh1542_wm36_12_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_c19(1);
   bh1542_wm35_11_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1796: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1796_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_copy1797_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1796_Out0_copy1797_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1798_In0_c20 <= "" & bh1542_wm36_0_c20 & bh1542_wm36_1_c20 & bh1542_wm36_2_c20 & bh1542_wm36_3_c20 & bh1542_wm36_4_c20 & bh1542_wm36_5_c20;
   bh1542_wm36_13_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_c20(0);
   bh1542_wm35_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_c20(1);
   bh1542_wm34_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1798: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1798_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_copy1799_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1798_Out0_copy1799_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In0_c19 <= "" & bh1542_wm36_6_c19 & bh1542_wm36_7_c19 & bh1542_wm36_8_c19 & bh1542_wm36_9_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In1_c20 <= "" & bh1542_wm35_0_c20;
   bh1542_wm36_14_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_c20(0);
   bh1542_wm35_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_c20(1);
   bh1542_wm34_12_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1800: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1800_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_copy1801_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1800_Out0_copy1801_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1802_In0_c19 <= "" & bh1542_wm35_1_c19 & bh1542_wm35_2_c19 & bh1542_wm35_3_c19 & bh1542_wm35_4_c19 & bh1542_wm35_5_c19 & bh1542_wm35_6_c19;
   bh1542_wm35_14_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_c19(0);
   bh1542_wm34_13_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_c19(1);
   bh1542_wm33_12_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1802: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1802_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_copy1803_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1802_Out0_copy1803_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1804_In0_c19 <= "" & bh1542_wm35_7_c19 & bh1542_wm35_8_c19 & bh1542_wm35_9_c19;
   bh1542_wm35_15_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_c19(0);
   bh1542_wm34_14_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1804: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1804_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_copy1805_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1804_Out0_copy1805_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1806_In0_c20 <= "" & bh1542_wm34_0_c20 & bh1542_wm34_1_c20 & bh1542_wm34_2_c20 & bh1542_wm34_3_c20 & bh1542_wm34_4_c20 & bh1542_wm34_5_c20;
   bh1542_wm34_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_c20(0);
   bh1542_wm33_13_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_c20(1);
   bh1542_wm32_10_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1806: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1806_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_copy1807_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1806_Out0_copy1807_c20; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1809_bh1542_uid1810_In0_c19 <= "" & bh1542_wm34_6_c19 & bh1542_wm34_7_c19 & bh1542_wm34_8_c19 & bh1542_wm34_9_c19 & bh1542_wm34_10_c19;
   bh1542_wm34_16_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_c19(0);
   bh1542_wm33_14_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_c19(1);
   bh1542_wm32_11_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_c19(2);
   Compressor_5_3_Freq300_uid1809_uid1810: Compressor_5_3_Freq300_uid1809
      port map ( X0 => Compressor_5_3_Freq300_uid1809_bh1542_uid1810_In0_c19,
                 R => Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_copy1811_c19);
   Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1810_Out0_copy1811_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1812_In0_c20 <= "" & bh1542_wm33_0_c20 & bh1542_wm33_1_c20 & bh1542_wm33_2_c20 & bh1542_wm33_3_c20 & bh1542_wm33_4_c20 & bh1542_wm33_5_c20;
   bh1542_wm33_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_c20(0);
   bh1542_wm32_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_c20(1);
   bh1542_wm31_10_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1812: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1812_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_copy1813_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1812_Out0_copy1813_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1814_In0_c19 <= "" & bh1542_wm33_6_c19 & bh1542_wm33_7_c19 & bh1542_wm33_8_c19 & bh1542_wm33_9_c19 & bh1542_wm33_10_c19 & bh1542_wm33_11_c19;
   bh1542_wm33_16_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_c19(0);
   bh1542_wm32_13_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_c19(1);
   bh1542_wm31_11_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1814: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1814_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_copy1815_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1814_Out0_copy1815_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1816_In0_c20 <= "" & bh1542_wm32_0_c20 & bh1542_wm32_1_c20 & bh1542_wm32_2_c20 & bh1542_wm32_3_c20 & bh1542_wm32_4_c20 & bh1542_wm32_5_c20;
   bh1542_wm32_14_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_c20(0);
   bh1542_wm31_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_c20(1);
   bh1542_wm30_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1816: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1816_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_copy1817_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1816_Out0_copy1817_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In0_c19 <= "" & bh1542_wm32_6_c19 & bh1542_wm32_7_c19 & bh1542_wm32_8_c19 & bh1542_wm32_9_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In1_c20 <= "" & bh1542_wm31_0_c20;
   bh1542_wm32_15_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_c20(0);
   bh1542_wm31_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_c20(1);
   bh1542_wm30_12_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1818: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1818_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_copy1819_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1818_Out0_copy1819_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1820_In0_c19 <= "" & bh1542_wm31_1_c19 & bh1542_wm31_2_c19 & bh1542_wm31_3_c19 & bh1542_wm31_4_c19 & bh1542_wm31_5_c19 & bh1542_wm31_6_c19;
   bh1542_wm31_14_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_c19(0);
   bh1542_wm30_13_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_c19(1);
   bh1542_wm29_12_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1820: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1820_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_copy1821_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1820_Out0_copy1821_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1822_In0_c19 <= "" & bh1542_wm31_7_c19 & bh1542_wm31_8_c19 & bh1542_wm31_9_c19;
   bh1542_wm31_15_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_c19(0);
   bh1542_wm30_14_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1822: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1822_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_copy1823_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1822_Out0_copy1823_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1824_In0_c20 <= "" & bh1542_wm30_0_c20 & bh1542_wm30_1_c20 & bh1542_wm30_2_c20 & bh1542_wm30_3_c20 & bh1542_wm30_4_c20 & bh1542_wm30_5_c20;
   bh1542_wm30_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_c20(0);
   bh1542_wm29_13_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_c20(1);
   bh1542_wm28_10_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1824: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1824_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_copy1825_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1824_Out0_copy1825_c20; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1809_bh1542_uid1826_In0_c19 <= "" & bh1542_wm30_6_c19 & bh1542_wm30_7_c19 & bh1542_wm30_8_c19 & bh1542_wm30_9_c19 & bh1542_wm30_10_c19;
   bh1542_wm30_16_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_c19(0);
   bh1542_wm29_14_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_c19(1);
   bh1542_wm28_11_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_c19(2);
   Compressor_5_3_Freq300_uid1809_uid1826: Compressor_5_3_Freq300_uid1809
      port map ( X0 => Compressor_5_3_Freq300_uid1809_bh1542_uid1826_In0_c19,
                 R => Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_copy1827_c19);
   Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_c19 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1826_Out0_copy1827_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1828_In0_c20 <= "" & bh1542_wm29_0_c20 & bh1542_wm29_1_c20 & bh1542_wm29_2_c20 & bh1542_wm29_3_c20 & bh1542_wm29_4_c20 & bh1542_wm29_5_c20;
   bh1542_wm29_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_c20(0);
   bh1542_wm28_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_c20(1);
   bh1542_wm27_10_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1828: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1828_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_copy1829_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1828_Out0_copy1829_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1830_In0_c19 <= "" & bh1542_wm29_6_c19 & bh1542_wm29_7_c19 & bh1542_wm29_8_c19 & bh1542_wm29_9_c19 & bh1542_wm29_10_c19 & bh1542_wm29_11_c19;
   bh1542_wm29_16_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_c19(0);
   bh1542_wm28_13_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_c19(1);
   bh1542_wm27_11_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1830: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1830_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_copy1831_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1830_Out0_copy1831_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1832_In0_c20 <= "" & bh1542_wm28_0_c20 & bh1542_wm28_1_c20 & bh1542_wm28_2_c20 & bh1542_wm28_3_c20 & bh1542_wm28_4_c20 & bh1542_wm28_5_c20;
   bh1542_wm28_14_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_c20(0);
   bh1542_wm27_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_c20(1);
   bh1542_wm26_11_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1832: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1832_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_copy1833_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1832_Out0_copy1833_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In0_c19 <= "" & bh1542_wm28_6_c19 & bh1542_wm28_7_c19 & bh1542_wm28_8_c19 & bh1542_wm28_9_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In1_c20 <= "" & bh1542_wm27_0_c20;
   bh1542_wm28_15_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_c20(0);
   bh1542_wm27_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_c20(1);
   bh1542_wm26_12_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1834: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1834_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_copy1835_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1834_Out0_copy1835_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1836_In0_c19 <= "" & bh1542_wm27_1_c19 & bh1542_wm27_2_c19 & bh1542_wm27_3_c19 & bh1542_wm27_4_c19 & bh1542_wm27_5_c19 & bh1542_wm27_6_c19;
   bh1542_wm27_14_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_c19(0);
   bh1542_wm26_13_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_c19(1);
   bh1542_wm25_11_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1836: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1836_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_copy1837_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1836_Out0_copy1837_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1838_In0_c19 <= "" & bh1542_wm27_7_c19 & bh1542_wm27_8_c19 & bh1542_wm27_9_c19;
   bh1542_wm27_15_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_c19(0);
   bh1542_wm26_14_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1838: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1838_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_copy1839_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1838_Out0_copy1839_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1840_In0_c20 <= "" & bh1542_wm26_0_c20 & bh1542_wm26_1_c20 & bh1542_wm26_2_c20 & bh1542_wm26_3_c20 & bh1542_wm26_4_c20 & bh1542_wm26_5_c20;
   bh1542_wm26_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_c20(0);
   bh1542_wm25_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_c20(1);
   bh1542_wm24_8_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1840: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1840_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_copy1841_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1840_Out0_copy1841_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In0_c19 <= "" & bh1542_wm26_6_c19 & bh1542_wm26_7_c19 & bh1542_wm26_8_c19 & bh1542_wm26_9_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In1_c20 <= "" & bh1542_wm25_0_c20;
   bh1542_wm26_16_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_c20(0);
   bh1542_wm25_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_c20(1);
   bh1542_wm24_9_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1842: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1842_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_copy1843_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1842_Out0_copy1843_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1844_In0_c19 <= "" & bh1542_wm25_1_c19 & bh1542_wm25_2_c19 & bh1542_wm25_3_c19 & bh1542_wm25_4_c19 & bh1542_wm25_5_c19 & bh1542_wm25_6_c19;
   bh1542_wm25_14_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_c19(0);
   bh1542_wm24_10_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_c19(1);
   bh1542_wm23_8_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1844: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1844_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_copy1845_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1844_Out0_copy1845_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1846_In0_c19 <= "" & bh1542_wm25_7_c19 & bh1542_wm25_8_c19 & bh1542_wm25_9_c19 & bh1542_wm25_10_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1846_In1_c19 <= "" & bh1542_wm24_0_c19;
   bh1542_wm25_15_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_c19(0);
   bh1542_wm24_11_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_c19(1);
   bh1542_wm23_9_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1846: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1846_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1846_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_copy1847_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1846_Out0_copy1847_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1848_In0_c19 <= "" & bh1542_wm24_1_c19 & bh1542_wm24_2_c19 & bh1542_wm24_3_c19 & bh1542_wm24_4_c19 & bh1542_wm24_5_c19 & bh1542_wm24_6_c19;
   bh1542_wm24_12_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_c19(0);
   bh1542_wm23_10_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_c19(1);
   bh1542_wm22_8_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1848: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1848_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_copy1849_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1848_Out0_copy1849_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1850_In0_c19 <= "" & bh1542_wm23_0_c19 & bh1542_wm23_1_c19 & bh1542_wm23_2_c19 & bh1542_wm23_3_c19 & bh1542_wm23_4_c19 & "0";
   bh1542_wm23_11_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_c19(0);
   bh1542_wm22_9_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_c19(1);
   bh1542_wm21_6_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1850: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1850_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_copy1851_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1850_Out0_copy1851_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1852_In0_c19 <= "" & bh1542_wm23_5_c19 & bh1542_wm23_6_c19 & bh1542_wm23_7_c19;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1852_In1_c19 <= "" & bh1542_wm22_0_c19 & bh1542_wm22_1_c19;
   bh1542_wm23_12_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_c19(0);
   bh1542_wm22_10_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_c19(1);
   bh1542_wm21_7_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_c19(2);
   Compressor_23_3_Freq300_uid1759_uid1852: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1852_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1852_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_copy1853_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1852_Out0_copy1853_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1854_In0_c19 <= "" & bh1542_wm22_2_c19 & bh1542_wm22_3_c19 & bh1542_wm22_4_c19 & bh1542_wm22_5_c19 & bh1542_wm22_6_c19 & bh1542_wm22_7_c19;
   bh1542_wm22_11_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_c19(0);
   bh1542_wm21_8_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_c19(1);
   bh1542_wm20_6_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1854: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1854_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_copy1855_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1854_Out0_copy1855_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1856_In0_c19 <= "" & bh1542_wm21_0_c19 & bh1542_wm21_1_c19 & bh1542_wm21_2_c19 & bh1542_wm21_3_c19 & bh1542_wm21_4_c19 & bh1542_wm21_5_c19;
   bh1542_wm21_9_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_c19(0);
   bh1542_wm20_7_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_c19(1);
   bh1542_wm19_5_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1856: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1856_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_copy1857_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1856_Out0_copy1857_c19; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1858_In0_c19 <= "" & bh1542_wm20_0_c19 & bh1542_wm20_1_c19 & bh1542_wm20_2_c19 & bh1542_wm20_3_c19 & bh1542_wm20_4_c19 & bh1542_wm20_5_c19;
   bh1542_wm20_8_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_c19(0);
   bh1542_wm19_6_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_c19(1);
   bh1542_wm18_4_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_c19(2);
   Compressor_6_3_Freq300_uid1775_uid1858: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1858_In0_c19,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_copy1859_c19);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_c19 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1858_Out0_copy1859_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1860_In0_c19 <= "" & bh1542_wm19_0_c19 & bh1542_wm19_1_c19 & bh1542_wm19_2_c19 & bh1542_wm19_3_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1860_In1_c19 <= "" & bh1542_wm18_0_c19;
   bh1542_wm19_7_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_c19(0);
   bh1542_wm18_5_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_c19(1);
   bh1542_wm17_3_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1860: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1860_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1860_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_copy1861_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1860_Out0_copy1861_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1862_In0_c19 <= "" & bh1542_wm18_1_c19 & bh1542_wm18_2_c19 & bh1542_wm18_3_c19;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1862_In1_c19 <= "" & bh1542_wm17_0_c19 & bh1542_wm17_1_c19;
   bh1542_wm18_6_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_c19(0);
   bh1542_wm17_4_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_c19(1);
   bh1542_wm16_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_c19(2);
   Compressor_23_3_Freq300_uid1759_uid1862: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1862_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1862_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_copy1863_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1862_Out0_copy1863_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1864_In0_c19 <= "" & bh1542_wm16_0_c19 & bh1542_wm16_1_c19 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1864_In1_c19 <= "" & bh1542_wm15_0_c19 & bh1542_wm15_1_c19;
   bh1542_wm16_3_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_c19(0);
   bh1542_wm15_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_c19(1);
   bh1542_wm14_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_c19(2);
   Compressor_23_3_Freq300_uid1759_uid1864: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1864_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1864_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_copy1865_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1864_Out0_copy1865_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1866_In0_c19 <= "" & bh1542_wm14_0_c19 & bh1542_wm14_1_c19 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1866_In1_c19 <= "" & bh1542_wm13_0_c19 & bh1542_wm13_1_c19;
   bh1542_wm14_3_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_c19(0);
   bh1542_wm13_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_c19(1);
   bh1542_wm12_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_c19(2);
   Compressor_23_3_Freq300_uid1759_uid1866: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1866_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1866_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_copy1867_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1866_Out0_copy1867_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1868_In0_c19 <= "" & bh1542_wm12_0_c19 & bh1542_wm12_1_c19 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1868_In1_c19 <= "" & bh1542_wm11_0_c19 & bh1542_wm11_1_c19;
   bh1542_wm12_3_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_c19(0);
   bh1542_wm11_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_c19(1);
   bh1542_wm10_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_c19(2);
   Compressor_23_3_Freq300_uid1759_uid1868: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1868_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1868_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_copy1869_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1868_Out0_copy1869_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1870_In0_c19 <= "" & bh1542_wm10_0_c19 & bh1542_wm10_1_c19 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1870_In1_c19 <= "" & bh1542_wm9_0_c19 & bh1542_wm9_1_c19;
   bh1542_wm10_3_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_c19(0);
   bh1542_wm9_2_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_c19(1);
   Compressor_23_3_Freq300_uid1759_uid1870: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1870_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1870_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_copy1871_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1870_Out0_copy1871_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1872_In0_c20 <= "" & bh1542_wm46_3_c20 & bh1542_wm46_4_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1872_In1_c20 <= "" & bh1542_wm45_4_c20 & bh1542_wm45_5_c20;
   bh1542_wm46_5_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_c20(0);
   bh1542_wm45_6_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_c20(1);
   bh1542_wm44_7_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1872: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1872_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1872_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_copy1873_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1872_Out0_copy1873_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1874_In0_c20 <= "" & bh1542_wm44_5_c20 & bh1542_wm44_6_c20 & "0";
   bh1542_wm44_8_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_c20(0);
   bh1542_wm43_8_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1874: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1874_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_copy1875_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1874_Out0_copy1875_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1876_In0_c20 <= "" & bh1542_wm43_5_c20 & bh1542_wm43_6_c20 & bh1542_wm43_7_c20;
   bh1542_wm43_9_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_c20(0);
   bh1542_wm42_11_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1876: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1876_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_copy1877_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1876_Out0_copy1877_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1878_In0_c20 <= "" & bh1542_wm42_7_c20 & bh1542_wm42_8_c20 & bh1542_wm42_9_c20 & bh1542_wm42_10_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1878_In1_c20 <= "" & bh1542_wm41_9_c20;
   bh1542_wm42_12_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_c20(0);
   bh1542_wm41_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_c20(1);
   bh1542_wm40_15_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1878: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1878_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1878_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_copy1879_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1878_Out0_copy1879_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1880_In0_c20 <= "" & bh1542_wm41_10_c20 & bh1542_wm41_11_c20 & bh1542_wm41_12_c20;
   bh1542_wm41_14_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_c20(0);
   bh1542_wm40_16_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1880: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1880_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_copy1881_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1880_Out0_copy1881_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1882_In0_c20 <= "" & bh1542_wm40_10_c20 & bh1542_wm40_11_c20 & bh1542_wm40_12_c20 & bh1542_wm40_13_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1882_In1_c20 <= "" & bh1542_wm39_11_c20;
   bh1542_wm40_17_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_c20(0);
   bh1542_wm39_16_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_c20(1);
   bh1542_wm38_17_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1882: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1882_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1882_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_copy1883_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1882_Out0_copy1883_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In0_c20 <= "" & bh1542_wm39_12_c20 & bh1542_wm39_13_c20 & bh1542_wm39_14_c20 & bh1542_wm39_15_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In1_c19 <= "" & bh1542_wm38_16_c19;
   bh1542_wm39_17_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_c20(0);
   bh1542_wm38_18_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_c20(1);
   bh1542_wm37_18_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1884: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1884_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_copy1885_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1884_Out0_copy1885_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1886_In0_c20 <= "" & bh1542_wm38_15_c20 & bh1542_wm38_14_c20 & bh1542_wm38_13_c20 & bh1542_wm38_12_c20 & bh1542_wm38_11_c20 & bh1542_wm38_10_c20;
   bh1542_wm38_19_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_c20(0);
   bh1542_wm37_19_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_c20(1);
   bh1542_wm36_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1886: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1886_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_copy1887_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1886_Out0_copy1887_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1888_In0_c20 <= "" & bh1542_wm37_17_c20 & bh1542_wm37_12_c20 & bh1542_wm37_13_c20 & bh1542_wm37_14_c20 & bh1542_wm37_15_c20 & bh1542_wm37_16_c20;
   bh1542_wm37_20_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_c20(0);
   bh1542_wm36_16_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_c20(1);
   bh1542_wm35_16_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1888: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1888_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_copy1889_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1888_Out0_copy1889_c20; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1809_bh1542_uid1890_In0_c20 <= "" & bh1542_wm36_10_c20 & bh1542_wm36_11_c20 & bh1542_wm36_12_c20 & bh1542_wm36_13_c20 & bh1542_wm36_14_c20;
   bh1542_wm36_17_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_c20(0);
   bh1542_wm35_17_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_c20(1);
   bh1542_wm34_17_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_c20(2);
   Compressor_5_3_Freq300_uid1809_uid1890: Compressor_5_3_Freq300_uid1809
      port map ( X0 => Compressor_5_3_Freq300_uid1809_bh1542_uid1890_In0_c20,
                 R => Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_copy1891_c20);
   Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1890_Out0_copy1891_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1892_In0_c20 <= "" & bh1542_wm35_10_c20 & bh1542_wm35_11_c20 & bh1542_wm35_12_c20 & bh1542_wm35_13_c20 & bh1542_wm35_14_c20 & bh1542_wm35_15_c20;
   bh1542_wm35_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_c20(0);
   bh1542_wm34_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_c20(1);
   bh1542_wm33_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1892: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1892_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_copy1893_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1892_Out0_copy1893_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1894_In0_c20 <= "" & bh1542_wm34_16_c20 & bh1542_wm34_15_c20 & bh1542_wm34_14_c20 & bh1542_wm34_13_c20 & bh1542_wm34_12_c20 & bh1542_wm34_11_c20;
   bh1542_wm34_19_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_c20(0);
   bh1542_wm33_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_c20(1);
   bh1542_wm32_16_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1894: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1894_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_copy1895_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1894_Out0_copy1895_c20; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1809_bh1542_uid1896_In0_c20 <= "" & bh1542_wm33_16_c20 & bh1542_wm33_15_c20 & bh1542_wm33_14_c20 & bh1542_wm33_13_c20 & bh1542_wm33_12_c20;
   bh1542_wm33_19_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_c20(0);
   bh1542_wm32_17_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_c20(1);
   bh1542_wm31_16_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_c20(2);
   Compressor_5_3_Freq300_uid1809_uid1896: Compressor_5_3_Freq300_uid1809
      port map ( X0 => Compressor_5_3_Freq300_uid1809_bh1542_uid1896_In0_c20,
                 R => Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_copy1897_c20);
   Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1896_Out0_copy1897_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1898_In0_c20 <= "" & bh1542_wm32_10_c20 & bh1542_wm32_11_c20 & bh1542_wm32_12_c20 & bh1542_wm32_13_c20 & bh1542_wm32_14_c20 & bh1542_wm32_15_c20;
   bh1542_wm32_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_c20(0);
   bh1542_wm31_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_c20(1);
   bh1542_wm30_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1898: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1898_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_copy1899_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1898_Out0_copy1899_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1900_In0_c20 <= "" & bh1542_wm31_10_c20 & bh1542_wm31_11_c20 & bh1542_wm31_12_c20 & bh1542_wm31_13_c20 & bh1542_wm31_14_c20 & bh1542_wm31_15_c20;
   bh1542_wm31_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_c20(0);
   bh1542_wm30_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_c20(1);
   bh1542_wm29_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1900: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1900_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_copy1901_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1900_Out0_copy1901_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1902_In0_c20 <= "" & bh1542_wm30_16_c20 & bh1542_wm30_15_c20 & bh1542_wm30_14_c20 & bh1542_wm30_13_c20 & bh1542_wm30_12_c20 & bh1542_wm30_11_c20;
   bh1542_wm30_19_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_c20(0);
   bh1542_wm29_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_c20(1);
   bh1542_wm28_16_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1902: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1902_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_copy1903_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1902_Out0_copy1903_c20; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1809_bh1542_uid1904_In0_c20 <= "" & bh1542_wm29_16_c20 & bh1542_wm29_15_c20 & bh1542_wm29_14_c20 & bh1542_wm29_13_c20 & bh1542_wm29_12_c20;
   bh1542_wm29_19_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_c20(0);
   bh1542_wm28_17_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_c20(1);
   bh1542_wm27_16_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_c20(2);
   Compressor_5_3_Freq300_uid1809_uid1904: Compressor_5_3_Freq300_uid1809
      port map ( X0 => Compressor_5_3_Freq300_uid1809_bh1542_uid1904_In0_c20,
                 R => Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_copy1905_c20);
   Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1904_Out0_copy1905_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1906_In0_c20 <= "" & bh1542_wm28_10_c20 & bh1542_wm28_11_c20 & bh1542_wm28_12_c20 & bh1542_wm28_13_c20 & bh1542_wm28_14_c20 & bh1542_wm28_15_c20;
   bh1542_wm28_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_c20(0);
   bh1542_wm27_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_c20(1);
   bh1542_wm26_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1906: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1906_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_copy1907_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1906_Out0_copy1907_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1908_In0_c20 <= "" & bh1542_wm27_10_c20 & bh1542_wm27_11_c20 & bh1542_wm27_12_c20 & bh1542_wm27_13_c20 & bh1542_wm27_14_c20 & bh1542_wm27_15_c20;
   bh1542_wm27_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_c20(0);
   bh1542_wm26_18_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_c20(1);
   bh1542_wm25_16_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1908: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1908_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_copy1909_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1908_Out0_copy1909_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1910_In0_c20 <= "" & bh1542_wm26_16_c20 & bh1542_wm26_15_c20 & bh1542_wm26_14_c20 & bh1542_wm26_13_c20 & bh1542_wm26_12_c20 & bh1542_wm26_11_c20;
   bh1542_wm26_19_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_c20(0);
   bh1542_wm25_17_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_c20(1);
   bh1542_wm24_13_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1910: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1910_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_copy1911_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1910_Out0_copy1911_c20; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1809_bh1542_uid1912_In0_c20 <= "" & bh1542_wm25_11_c20 & bh1542_wm25_12_c20 & bh1542_wm25_13_c20 & bh1542_wm25_14_c20 & bh1542_wm25_15_c20;
   bh1542_wm25_18_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_c20(0);
   bh1542_wm24_14_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_c20(1);
   bh1542_wm23_13_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_c20(2);
   Compressor_5_3_Freq300_uid1809_uid1912: Compressor_5_3_Freq300_uid1809
      port map ( X0 => Compressor_5_3_Freq300_uid1809_bh1542_uid1912_In0_c20,
                 R => Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_copy1913_c20);
   Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_c20 <= Compressor_5_3_Freq300_uid1809_bh1542_uid1912_Out0_copy1913_c20; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1775_bh1542_uid1914_In0_c20 <= "" & bh1542_wm24_7_c20 & bh1542_wm24_8_c20 & bh1542_wm24_9_c20 & bh1542_wm24_10_c20 & bh1542_wm24_11_c20 & bh1542_wm24_12_c20;
   bh1542_wm24_15_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_c20(0);
   bh1542_wm23_14_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_c20(1);
   bh1542_wm22_12_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_c20(2);
   Compressor_6_3_Freq300_uid1775_uid1914: Compressor_6_3_Freq300_uid1775
      port map ( X0 => Compressor_6_3_Freq300_uid1775_bh1542_uid1914_In0_c20,
                 R => Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_copy1915_c20);
   Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_c20 <= Compressor_6_3_Freq300_uid1775_bh1542_uid1914_Out0_copy1915_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1916_In0_c19 <= "" & bh1542_wm23_8_c19 & bh1542_wm23_9_c19 & bh1542_wm23_10_c19 & bh1542_wm23_11_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1916_In1_c19 <= "" & bh1542_wm22_8_c19;
   bh1542_wm23_15_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_c19(0);
   bh1542_wm22_13_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_c19(1);
   bh1542_wm21_10_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1916: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1916_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1916_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_copy1917_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1916_Out0_copy1917_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1918_In0_c19 <= "" & bh1542_wm22_9_c19 & bh1542_wm22_10_c19 & bh1542_wm22_11_c19;
   bh1542_wm22_14_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_c19(0);
   bh1542_wm21_11_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1918: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1918_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_copy1919_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1918_Out0_copy1919_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In0_c19 <= "" & bh1542_wm21_6_c19 & bh1542_wm21_7_c19 & bh1542_wm21_8_c19 & bh1542_wm21_9_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c0 <= "" & "0";
   bh1542_wm21_12_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_c19(0);
   bh1542_wm20_9_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_c19(1);
   bh1542_wm19_8_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1920: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1920_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_copy1921_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1920_Out0_copy1921_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1922_In0_c19 <= "" & bh1542_wm20_6_c19 & bh1542_wm20_7_c19 & bh1542_wm20_8_c19;
   bh1542_wm20_10_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_c19(0);
   bh1542_wm19_9_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1922: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1922_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_copy1923_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1922_Out0_copy1923_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In0_c19 <= "" & bh1542_wm19_4_c19 & bh1542_wm19_5_c19 & bh1542_wm19_6_c19 & bh1542_wm19_7_c19;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c0 <= "" & "0";
   bh1542_wm19_10_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_c19(0);
   bh1542_wm18_7_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_c19(1);
   bh1542_wm17_5_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1924: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1924_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_copy1925_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1924_Out0_copy1925_c19; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1926_In0_c19 <= "" & bh1542_wm18_4_c19 & bh1542_wm18_5_c19 & bh1542_wm18_6_c19;
   bh1542_wm18_8_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_c19(0);
   bh1542_wm17_6_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_c19(1);
   Compressor_3_2_Freq300_uid1763_uid1926: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1926_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_copy1927_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_c19 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1926_Out0_copy1927_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1928_In0_c19 <= "" & bh1542_wm17_2_c19 & bh1542_wm17_3_c19 & bh1542_wm17_4_c19;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1928_In1_c19 <= "" & bh1542_wm16_2_c19 & bh1542_wm16_3_c19;
   bh1542_wm17_7_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_c19(0);
   bh1542_wm16_4_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_c19(1);
   bh1542_wm15_3_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_c19(2);
   Compressor_23_3_Freq300_uid1759_uid1928: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1928_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1928_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_copy1929_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_c19 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1928_Out0_copy1929_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1930_In0_c19 <= "" & bh1542_wm14_2_c19 & bh1542_wm14_3_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1930_In1_c19 <= "" & bh1542_wm13_2_c19;
   bh1542_wm14_4_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_c19(0);
   bh1542_wm13_3_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_c19(1);
   bh1542_wm12_4_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1930: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1930_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1930_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_copy1931_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1930_Out0_copy1931_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1932_In0_c19 <= "" & bh1542_wm12_2_c19 & bh1542_wm12_3_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1932_In1_c19 <= "" & bh1542_wm11_2_c19;
   bh1542_wm12_5_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_c19(0);
   bh1542_wm11_3_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_c19(1);
   bh1542_wm10_4_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_c19(2);
   Compressor_14_3_Freq300_uid1767_uid1932: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1932_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1932_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_copy1933_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1932_Out0_copy1933_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1934_In0_c19 <= "" & bh1542_wm10_2_c19 & bh1542_wm10_3_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1934_In1_c19 <= "" & bh1542_wm9_2_c19;
   bh1542_wm10_5_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_c19(0);
   bh1542_wm9_3_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_c19(1);
   Compressor_14_3_Freq300_uid1767_uid1934: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1934_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1934_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_copy1935_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1934_Out0_copy1935_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1936_In0_c20 <= "" & bh1542_wm44_7_c20 & bh1542_wm44_8_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1936_In1_c20 <= "" & bh1542_wm43_8_c20 & bh1542_wm43_9_c20;
   bh1542_wm44_9_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_c20(0);
   bh1542_wm43_10_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_c20(1);
   bh1542_wm42_13_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1936: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1936_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1936_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_copy1937_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1936_Out0_copy1937_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1938_In0_c20 <= "" & bh1542_wm42_11_c20 & bh1542_wm42_12_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1938_In1_c20 <= "" & bh1542_wm41_13_c20 & bh1542_wm41_14_c20;
   bh1542_wm42_14_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_c20(0);
   bh1542_wm41_15_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_c20(1);
   bh1542_wm40_18_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1938: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1938_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1938_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_copy1939_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1938_Out0_copy1939_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1940_In0_c20 <= "" & bh1542_wm40_14_c20 & bh1542_wm40_15_c20 & bh1542_wm40_16_c20 & bh1542_wm40_17_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1940_In1_c20 <= "" & bh1542_wm39_16_c20;
   bh1542_wm40_19_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_c20(0);
   bh1542_wm39_18_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_c20(1);
   bh1542_wm38_20_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1940: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1940_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1940_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_copy1941_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1940_Out0_copy1941_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1942_In0_c20 <= "" & bh1542_wm38_17_c20 & bh1542_wm38_18_c20 & bh1542_wm38_19_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1942_In1_c20 <= "" & bh1542_wm37_18_c20 & bh1542_wm37_19_c20;
   bh1542_wm38_21_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_c20(0);
   bh1542_wm37_21_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_c20(1);
   bh1542_wm36_18_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1942: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1942_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1942_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_copy1943_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1942_Out0_copy1943_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1944_In0_c20 <= "" & bh1542_wm36_15_c20 & bh1542_wm36_16_c20 & bh1542_wm36_17_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1944_In1_c20 <= "" & bh1542_wm35_16_c20 & bh1542_wm35_17_c20;
   bh1542_wm36_19_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_c20(0);
   bh1542_wm35_19_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_c20(1);
   bh1542_wm34_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1944: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1944_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1944_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_copy1945_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1944_Out0_copy1945_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1946_In0_c20 <= "" & bh1542_wm34_17_c20 & bh1542_wm34_18_c20 & bh1542_wm34_19_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1946_In1_c20 <= "" & bh1542_wm33_17_c20 & bh1542_wm33_18_c20;
   bh1542_wm34_21_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_c20(0);
   bh1542_wm33_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_c20(1);
   bh1542_wm32_19_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1946: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1946_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1946_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_copy1947_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1946_Out0_copy1947_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1948_In0_c20 <= "" & bh1542_wm32_16_c20 & bh1542_wm32_17_c20 & bh1542_wm32_18_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1948_In1_c20 <= "" & bh1542_wm31_16_c20 & bh1542_wm31_17_c20;
   bh1542_wm32_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_c20(0);
   bh1542_wm31_19_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_c20(1);
   bh1542_wm30_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1948: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1948_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1948_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_copy1949_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1948_Out0_copy1949_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1950_In0_c20 <= "" & bh1542_wm30_17_c20 & bh1542_wm30_18_c20 & bh1542_wm30_19_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1950_In1_c20 <= "" & bh1542_wm29_17_c20 & bh1542_wm29_18_c20;
   bh1542_wm30_21_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_c20(0);
   bh1542_wm29_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_c20(1);
   bh1542_wm28_19_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1950: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1950_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1950_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_copy1951_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1950_Out0_copy1951_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1952_In0_c20 <= "" & bh1542_wm28_16_c20 & bh1542_wm28_17_c20 & bh1542_wm28_18_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1952_In1_c20 <= "" & bh1542_wm27_16_c20 & bh1542_wm27_17_c20;
   bh1542_wm28_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_c20(0);
   bh1542_wm27_19_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_c20(1);
   bh1542_wm26_20_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1952: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1952_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1952_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_copy1953_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1952_Out0_copy1953_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In0_c20 <= "" & bh1542_wm26_10_c20 & bh1542_wm26_17_c20 & bh1542_wm26_18_c20 & bh1542_wm26_19_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c0 <= "" & "0";
   bh1542_wm26_21_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_c20(0);
   bh1542_wm25_19_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_c20(1);
   bh1542_wm24_16_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1954: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1954_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_copy1955_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1954_Out0_copy1955_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1956_In0_c20 <= "" & bh1542_wm25_16_c20 & bh1542_wm25_17_c20 & bh1542_wm25_18_c20;
   bh1542_wm25_20_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_c20(0);
   bh1542_wm24_17_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1956: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1956_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_copy1957_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1956_Out0_copy1957_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1958_In0_c20 <= "" & bh1542_wm24_13_c20 & bh1542_wm24_14_c20 & bh1542_wm24_15_c20;
   bh1542_wm24_18_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_c20(0);
   bh1542_wm23_16_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1958: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1958_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_copy1959_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1958_Out0_copy1959_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In0_c20 <= "" & bh1542_wm23_12_c20 & bh1542_wm23_13_c20 & bh1542_wm23_14_c20 & bh1542_wm23_15_c20;
   Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c0 <= "" & "0";
   bh1542_wm23_17_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_c20(0);
   bh1542_wm22_15_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_c20(1);
   bh1542_wm21_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1960: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1960_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_copy1961_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1960_Out0_copy1961_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1962_In0_c20 <= "" & bh1542_wm22_12_c20 & bh1542_wm22_13_c20 & bh1542_wm22_14_c20;
   bh1542_wm22_16_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_c20(0);
   bh1542_wm21_14_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1962: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1962_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_copy1963_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1962_Out0_copy1963_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1964_In0_c19 <= "" & bh1542_wm21_10_c19 & bh1542_wm21_11_c19 & bh1542_wm21_12_c19;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1964_In1_c19 <= "" & bh1542_wm20_9_c19 & bh1542_wm20_10_c19;
   bh1542_wm21_15_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_c20(0);
   bh1542_wm20_11_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_c20(1);
   bh1542_wm19_11_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1964: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1964_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1964_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_copy1965_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1964_Out0_copy1965_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1966_In0_c19 <= "" & bh1542_wm19_8_c19 & bh1542_wm19_9_c19 & bh1542_wm19_10_c19;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1966_In1_c19 <= "" & bh1542_wm18_7_c19 & bh1542_wm18_8_c19;
   bh1542_wm19_12_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_c20(0);
   bh1542_wm18_9_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_c20(1);
   bh1542_wm17_8_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid1966: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1966_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1966_In1_c19,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_copy1967_c19);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1966_Out0_copy1967_c20; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1968_In0_c19 <= "" & bh1542_wm17_5_c19 & bh1542_wm17_6_c19 & bh1542_wm17_7_c19;
   bh1542_wm17_9_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_c20(0);
   bh1542_wm16_5_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_c20(1);
   Compressor_3_2_Freq300_uid1763_uid1968: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1968_In0_c19,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_copy1969_c19);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_c20 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1968_Out0_copy1969_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1970_In0_c19 <= "" & bh1542_wm15_2_c19 & bh1542_wm15_3_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1970_In1_c19 <= "" & bh1542_wm14_4_c19;
   bh1542_wm15_4_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_c20(0);
   bh1542_wm14_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_c20(1);
   bh1542_wm13_4_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1970: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1970_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1970_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_copy1971_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1970_Out0_copy1971_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1972_In0_c19 <= "" & bh1542_wm12_4_c19 & bh1542_wm12_5_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1972_In1_c19 <= "" & bh1542_wm11_3_c19;
   bh1542_wm12_6_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_c20(0);
   bh1542_wm11_4_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_c20(1);
   bh1542_wm10_6_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid1972: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1972_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1972_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_copy1973_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1972_Out0_copy1973_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1974_In0_c19 <= "" & bh1542_wm10_4_c19 & bh1542_wm10_5_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1974_In1_c19 <= "" & bh1542_wm9_3_c19;
   bh1542_wm10_7_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_c19(0);
   bh1542_wm9_4_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_c19(1);
   Compressor_14_3_Freq300_uid1767_uid1974: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1974_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1974_In1_c19,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_copy1975_c19);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_c19 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1974_Out0_copy1975_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid1976_In0_c20 <= "" & bh1542_wm42_13_c20 & bh1542_wm42_14_c20 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid1976_In1_c20 <= "" & bh1542_wm41_15_c20;
   bh1542_wm42_15_c21 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_c21(0);
   bh1542_wm41_16_c21 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_c21(1);
   bh1542_wm40_20_c21 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_c21(2);
   Compressor_14_3_Freq300_uid1767_uid1976: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid1976_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid1976_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_copy1977_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_c21 <= Compressor_14_3_Freq300_uid1767_bh1542_uid1976_Out0_copy1977_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1978_In0_c20 <= "" & bh1542_wm40_18_c20 & bh1542_wm40_19_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1978_In1_c20 <= "" & bh1542_wm39_17_c20 & bh1542_wm39_18_c20;
   bh1542_wm40_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_c21(0);
   bh1542_wm39_19_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_c21(1);
   bh1542_wm38_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1978: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1978_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1978_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_copy1979_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1978_Out0_copy1979_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1980_In0_c20 <= "" & bh1542_wm38_20_c20 & bh1542_wm38_21_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1980_In1_c20 <= "" & bh1542_wm37_20_c20 & bh1542_wm37_21_c20;
   bh1542_wm38_23_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_c21(0);
   bh1542_wm37_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_c21(1);
   bh1542_wm36_20_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1980: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1980_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1980_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_copy1981_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1980_Out0_copy1981_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1982_In0_c20 <= "" & bh1542_wm36_18_c20 & bh1542_wm36_19_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1982_In1_c20 <= "" & bh1542_wm35_18_c20 & bh1542_wm35_19_c20;
   bh1542_wm36_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_c21(0);
   bh1542_wm35_20_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_c21(1);
   bh1542_wm34_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1982: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1982_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1982_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_copy1983_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1982_Out0_copy1983_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1984_In0_c20 <= "" & bh1542_wm34_20_c20 & bh1542_wm34_21_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1984_In1_c20 <= "" & bh1542_wm33_19_c20 & bh1542_wm33_20_c20;
   bh1542_wm34_23_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_c21(0);
   bh1542_wm33_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_c21(1);
   bh1542_wm32_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1984: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1984_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1984_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_copy1985_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1984_Out0_copy1985_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1986_In0_c20 <= "" & bh1542_wm32_19_c20 & bh1542_wm32_20_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1986_In1_c20 <= "" & bh1542_wm31_18_c20 & bh1542_wm31_19_c20;
   bh1542_wm32_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_c21(0);
   bh1542_wm31_20_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_c21(1);
   bh1542_wm30_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1986: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1986_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1986_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_copy1987_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1986_Out0_copy1987_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1988_In0_c20 <= "" & bh1542_wm30_20_c20 & bh1542_wm30_21_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1988_In1_c20 <= "" & bh1542_wm29_19_c20 & bh1542_wm29_20_c20;
   bh1542_wm30_23_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_c21(0);
   bh1542_wm29_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_c21(1);
   bh1542_wm28_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1988: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1988_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1988_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_copy1989_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1988_Out0_copy1989_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1990_In0_c20 <= "" & bh1542_wm28_19_c20 & bh1542_wm28_20_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1990_In1_c20 <= "" & bh1542_wm27_18_c20 & bh1542_wm27_19_c20;
   bh1542_wm28_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_c21(0);
   bh1542_wm27_20_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_c21(1);
   bh1542_wm26_22_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1990: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1990_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1990_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_copy1991_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1990_Out0_copy1991_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1992_In0_c20 <= "" & bh1542_wm26_20_c20 & bh1542_wm26_21_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid1992_In1_c20 <= "" & bh1542_wm25_19_c20 & bh1542_wm25_20_c20;
   bh1542_wm26_23_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_c21(0);
   bh1542_wm25_21_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_c21(1);
   bh1542_wm24_19_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1992: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1992_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1992_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_copy1993_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1992_Out0_copy1993_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid1994_In0_c20 <= "" & bh1542_wm24_16_c20 & bh1542_wm24_17_c20 & bh1542_wm24_18_c20;
   Compressor_23_3_Freq300_uid1759_bh1542_uid1994_In1_c20 <= "" & bh1542_wm23_16_c20 & bh1542_wm23_17_c20;
   bh1542_wm24_20_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_c21(0);
   bh1542_wm23_18_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_c21(1);
   bh1542_wm22_17_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_c21(2);
   Compressor_23_3_Freq300_uid1759_uid1994: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid1994_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid1994_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_copy1995_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_c21 <= Compressor_23_3_Freq300_uid1759_bh1542_uid1994_Out0_copy1995_c21; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1996_In0_c20 <= "" & bh1542_wm22_15_c20 & bh1542_wm22_16_c20 & "0";
   bh1542_wm22_18_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_c21(0);
   bh1542_wm21_16_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_c21(1);
   Compressor_3_2_Freq300_uid1763_uid1996: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1996_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_copy1997_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1996_Out0_copy1997_c21; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1763_bh1542_uid1998_In0_c20 <= "" & bh1542_wm21_13_c20 & bh1542_wm21_14_c20 & bh1542_wm21_15_c20;
   bh1542_wm21_17_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_c21(0);
   bh1542_wm20_12_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_c21(1);
   Compressor_3_2_Freq300_uid1763_uid1998: Compressor_3_2_Freq300_uid1763
      port map ( X0 => Compressor_3_2_Freq300_uid1763_bh1542_uid1998_In0_c20,
                 R => Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_copy1999_c20);
   Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_c21 <= Compressor_3_2_Freq300_uid1763_bh1542_uid1998_Out0_copy1999_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid2000_In0_c20 <= "" & bh1542_wm19_11_c20 & bh1542_wm19_12_c20 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid2000_In1_c20 <= "" & bh1542_wm18_9_c20;
   bh1542_wm19_13_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_c20(0);
   bh1542_wm18_10_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_c20(1);
   bh1542_wm17_10_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid2000: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid2000_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid2000_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_copy2001_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2000_Out0_copy2001_c20; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1759_bh1542_uid2002_In0_c20 <= "" & bh1542_wm17_8_c20 & bh1542_wm17_9_c20 & "0";
   Compressor_23_3_Freq300_uid1759_bh1542_uid2002_In1_c20 <= "" & bh1542_wm16_4_c20 & bh1542_wm16_5_c20;
   bh1542_wm17_11_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_c20(0);
   bh1542_wm16_6_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_c20(1);
   bh1542_wm15_5_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_c20(2);
   Compressor_23_3_Freq300_uid1759_uid2002: Compressor_23_3_Freq300_uid1759
      port map ( X0 => Compressor_23_3_Freq300_uid1759_bh1542_uid2002_In0_c20,
                 X1 => Compressor_23_3_Freq300_uid1759_bh1542_uid2002_In1_c20,
                 R => Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_copy2003_c20);
   Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_c20 <= Compressor_23_3_Freq300_uid1759_bh1542_uid2002_Out0_copy2003_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid2004_In0_c20 <= "" & bh1542_wm13_3_c20 & bh1542_wm13_4_c20 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid2004_In1_c20 <= "" & bh1542_wm12_6_c20;
   bh1542_wm13_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_c20(0);
   bh1542_wm12_7_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_c20(1);
   bh1542_wm11_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_c20(2);
   Compressor_14_3_Freq300_uid1767_uid2004: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid2004_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid2004_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_copy2005_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2004_Out0_copy2005_c20; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In0_c20 <= "" & bh1542_wm10_6_c20 & bh1542_wm10_7_c20 & "0" & "0";
   Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In1_c19 <= "" & bh1542_wm9_4_c19;
   bh1542_wm10_8_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_c20(0);
   bh1542_wm9_5_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_c20(1);
   Compressor_14_3_Freq300_uid1767_uid2006: Compressor_14_3_Freq300_uid1767
      port map ( X0 => Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In0_c20,
                 X1 => Compressor_14_3_Freq300_uid1767_bh1542_uid2006_In1_c20,
                 R => Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_copy2007_c20);
   Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_c20 <= Compressor_14_3_Freq300_uid1767_bh1542_uid2006_Out0_copy2007_c20; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh1542_24_c21 <= bh1542_wm41_16_c21 & bh1542_wm42_15_c21 & bh1542_wm43_10_c21 & bh1542_wm44_9_c21 & bh1542_wm45_6_c21 & bh1542_wm46_5_c21 & bh1542_wm47_2_c21 & bh1542_wm48_2_c21 & bh1542_wm49_0_c21 & bh1542_wm50_0_c21 & bh1542_wm51_0_c21 & bh1542_wm52_0_c21 & bh1542_wm53_0_c21 & bh1542_wm54_0_c21 & bh1542_wm55_0_c21 & bh1542_wm56_0_c21 & bh1542_wm57_0_c21 & bh1542_wm58_0_c21 & bh1542_wm59_0_c21 & bh1542_wm60_0_c21 & bh1542_wm61_0_c21 & bh1542_wm62_0_c21 & bh1542_wm63_0_c21 & bh1542_wm64_0_c21 & bh1542_wm65_0_c21;

   bitheapFinalAdd_bh1542_In0_c21 <= "0" & bh1542_wm9_5_c21 & bh1542_wm10_8_c21 & bh1542_wm11_4_c21 & bh1542_wm12_7_c21 & bh1542_wm13_5_c21 & bh1542_wm14_5_c21 & bh1542_wm15_4_c21 & bh1542_wm16_6_c21 & bh1542_wm17_10_c21 & bh1542_wm18_10_c21 & bh1542_wm19_13_c21 & bh1542_wm20_11_c21 & bh1542_wm21_16_c21 & bh1542_wm22_17_c21 & bh1542_wm23_18_c21 & bh1542_wm24_19_c21 & bh1542_wm25_21_c21 & bh1542_wm26_22_c21 & bh1542_wm27_20_c21 & bh1542_wm28_21_c21 & bh1542_wm29_21_c21 & bh1542_wm30_22_c21 & bh1542_wm31_20_c21 & bh1542_wm32_21_c21 & bh1542_wm33_21_c21 & bh1542_wm34_22_c21 & bh1542_wm35_20_c21 & bh1542_wm36_20_c21 & bh1542_wm37_22_c21 & bh1542_wm38_22_c21 & bh1542_wm39_19_c21 & bh1542_wm40_20_c21;
   bitheapFinalAdd_bh1542_In1_c21 <= "0" & "0" & "0" & bh1542_wm11_5_c21 & "0" & "0" & "0" & bh1542_wm15_5_c21 & "0" & bh1542_wm17_11_c21 & "0" & "0" & bh1542_wm20_12_c21 & bh1542_wm21_17_c21 & bh1542_wm22_18_c21 & "0" & bh1542_wm24_20_c21 & "0" & bh1542_wm26_23_c21 & "0" & bh1542_wm28_22_c21 & "0" & bh1542_wm30_23_c21 & "0" & bh1542_wm32_22_c21 & "0" & bh1542_wm34_23_c21 & "0" & bh1542_wm36_21_c21 & "0" & bh1542_wm38_23_c21 & "0" & bh1542_wm40_21_c21;
   bitheapFinalAdd_bh1542_Cin_c0 <= '0';

   bitheapFinalAdd_bh1542: IntAdder_33_Freq300_uid2009
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 Cin => bitheapFinalAdd_bh1542_Cin_c0,
                 X => bitheapFinalAdd_bh1542_In0_c21,
                 Y => bitheapFinalAdd_bh1542_In1_c21,
                 R => bitheapFinalAdd_bh1542_Out_c21);
   bitheapResult_bh1542_c21 <= bitheapFinalAdd_bh1542_Out_c21(31 downto 0) & tmp_bitheapResult_bh1542_24_c21;
   RR_c21 <= signed(bitheapResult_bh1542_c21(56 downto 24));
R <= std_logic_vector(RR_c21);  
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid2014
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid2014 is
    port (clk, ce_20, ce_21, ce_22 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid2014 is
signal Mfull_c21, Mfull_c22 :  std_logic_vector(40 downto 0);
signal M_c22 :  std_logic_vector(40 downto 0);
signal X_c20, X_c21 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
            if ce_22 = '1' then
               Mfull_c22 <= Mfull_c21;
            end if;
         end if;
      end process;
   Mfull_c21 <= std_logic_vector(unsigned(X_c21) * unsigned(Y)); -- multiplier
   M_c22 <= Mfull_c22(40 downto 0);
   R <= M_c22;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_12x24_Freq300_uid2016
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_12x24_Freq300_uid2016 is
    port (clk, ce_20, ce_21, ce_22 : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of DSPBlock_12x24_Freq300_uid2016 is
signal Mfull_c21, Mfull_c22 :  std_logic_vector(36 downto 0);
signal M_c22 :  std_logic_vector(35 downto 0);
signal X_c20, X_c21 :  std_logic_vector(11 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
            if ce_22 = '1' then
               Mfull_c22 <= Mfull_c21;
            end if;
         end if;
      end process;
   Mfull_c21 <= std_logic_vector(signed(X_c21) * signed('0' & Y)); -- multiplier
   M_c22 <= Mfull_c22(35 downto 0);
   R <= M_c22;
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_1x1_signed_Freq300_uid2018
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_signed_Freq300_uid2018 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_signed_Freq300_uid2018 is
signal replicated_c19, replicated_c20, replicated_c21 :  std_logic_vector(0 downto 0);
signal prod_c21 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               replicated_c20 <= replicated_c19;
            end if;
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
         end if;
      end process;
   replicated_c19 <= (0 downto 0 => X(0));
   prod_c21 <= Y and replicated_c21;
   R <= prod_c21;
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid2020
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid2020 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid2020 is
   component MultTable_Freq300_uid2022 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2023_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2022
      port map ( X => Xtable_c21,
                 Y => Y1_copy2023_c21);
   Y1_c21 <= Y1_copy2023_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid2025
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid2025 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid2025 is
   component MultTable_Freq300_uid2027 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2028_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2027
      port map ( X => Xtable_c21,
                 Y => Y1_copy2028_c21);
   Y1_c21 <= Y1_copy2028_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid2030
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid2030 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid2030 is
   component MultTable_Freq300_uid2032 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2033_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2032
      port map ( X => Xtable_c21,
                 Y => Y1_copy2033_c21);
   Y1_c21 <= Y1_copy2033_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid2035
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid2035 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid2035 is
   component MultTable_Freq300_uid2037 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2038_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2037
      port map ( X => Xtable_c21,
                 Y => Y1_copy2038_c21);
   Y1_c21 <= Y1_copy2038_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2040
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2040 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2040 is
   component MultTable_Freq300_uid2042 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(3 downto 0);
signal Y1_c21 :  std_logic_vector(3 downto 0);
signal Y1_copy2043_c21 :  std_logic_vector(3 downto 0);
signal X_c20, X_c21 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2042
      port map ( X => Xtable_c21,
                 Y => Y1_copy2043_c21);
   Y1_c21 <= Y1_copy2043_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2045
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2045 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2045 is
   component MultTable_Freq300_uid2047 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2048_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2047
      port map ( X => Xtable_c21,
                 Y => Y1_copy2048_c21);
   Y1_c21 <= Y1_copy2048_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2050
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2050 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2050 is
   component MultTable_Freq300_uid2052 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2053_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2052
      port map ( X => Xtable_c21,
                 Y => Y1_copy2053_c21);
   Y1_c21 <= Y1_copy2053_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2055
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2055 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2055 is
   component MultTable_Freq300_uid2057 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2058_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2057
      port map ( X => Xtable_c21,
                 Y => Y1_copy2058_c21);
   Y1_c21 <= Y1_copy2058_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2060
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2060 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2060 is
   component MultTable_Freq300_uid2062 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2063_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2062
      port map ( X => Xtable_c21,
                 Y => Y1_copy2063_c21);
   Y1_c21 <= Y1_copy2063_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2065
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2065 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2065 is
   component MultTable_Freq300_uid2067 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2068_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2067
      port map ( X => Xtable_c21,
                 Y => Y1_copy2068_c21);
   Y1_c21 <= Y1_copy2068_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2070
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2070 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2070 is
   component MultTable_Freq300_uid2072 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(3 downto 0);
signal Y1_c21 :  std_logic_vector(3 downto 0);
signal Y1_copy2073_c21 :  std_logic_vector(3 downto 0);
signal X_c20, X_c21 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2072
      port map ( X => Xtable_c21,
                 Y => Y1_copy2073_c21);
   Y1_c21 <= Y1_copy2073_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2075
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2075 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2075 is
   component MultTable_Freq300_uid2077 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2078_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2077
      port map ( X => Xtable_c21,
                 Y => Y1_copy2078_c21);
   Y1_c21 <= Y1_copy2078_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2080
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2080 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2080 is
   component MultTable_Freq300_uid2082 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2083_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2082
      port map ( X => Xtable_c21,
                 Y => Y1_copy2083_c21);
   Y1_c21 <= Y1_copy2083_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2085
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2085 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2085 is
   component MultTable_Freq300_uid2087 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2088_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2087
      port map ( X => Xtable_c21,
                 Y => Y1_copy2088_c21);
   Y1_c21 <= Y1_copy2088_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2090
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2090 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2090 is
   component MultTable_Freq300_uid2092 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2093_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2092
      port map ( X => Xtable_c21,
                 Y => Y1_copy2093_c21);
   Y1_c21 <= Y1_copy2093_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2095
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2095 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2095 is
   component MultTable_Freq300_uid2097 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2098_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2097
      port map ( X => Xtable_c21,
                 Y => Y1_copy2098_c21);
   Y1_c21 <= Y1_copy2098_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2100
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2100 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2100 is
   component MultTable_Freq300_uid2102 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(3 downto 0);
signal Y1_c21 :  std_logic_vector(3 downto 0);
signal Y1_copy2103_c21 :  std_logic_vector(3 downto 0);
signal X_c20, X_c21 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2102
      port map ( X => Xtable_c21,
                 Y => Y1_copy2103_c21);
   Y1_c21 <= Y1_copy2103_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2105
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2105 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2105 is
   component MultTable_Freq300_uid2107 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2108_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2107
      port map ( X => Xtable_c21,
                 Y => Y1_copy2108_c21);
   Y1_c21 <= Y1_copy2108_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2110
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2110 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2110 is
   component MultTable_Freq300_uid2112 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2113_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2112
      port map ( X => Xtable_c21,
                 Y => Y1_copy2113_c21);
   Y1_c21 <= Y1_copy2113_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2115
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2115 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2115 is
   component MultTable_Freq300_uid2117 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2118_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2117
      port map ( X => Xtable_c21,
                 Y => Y1_copy2118_c21);
   Y1_c21 <= Y1_copy2118_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2120
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2120 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2120 is
   component MultTable_Freq300_uid2122 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2123_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2122
      port map ( X => Xtable_c21,
                 Y => Y1_copy2123_c21);
   Y1_c21 <= Y1_copy2123_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2125
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2125 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2125 is
   component MultTable_Freq300_uid2127 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2128_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2127
      port map ( X => Xtable_c21,
                 Y => Y1_copy2128_c21);
   Y1_c21 <= Y1_copy2128_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2130
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2130 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2130 is
   component MultTable_Freq300_uid2132 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(3 downto 0);
signal Y1_c21 :  std_logic_vector(3 downto 0);
signal Y1_copy2133_c21 :  std_logic_vector(3 downto 0);
signal X_c20, X_c21 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2132
      port map ( X => Xtable_c21,
                 Y => Y1_copy2133_c21);
   Y1_c21 <= Y1_copy2133_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2135
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2135 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2135 is
   component MultTable_Freq300_uid2137 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2138_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2137
      port map ( X => Xtable_c21,
                 Y => Y1_copy2138_c21);
   Y1_c21 <= Y1_copy2138_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2140
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2140 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2140 is
   component MultTable_Freq300_uid2142 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2143_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2142
      port map ( X => Xtable_c21,
                 Y => Y1_copy2143_c21);
   Y1_c21 <= Y1_copy2143_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2145
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2145 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2145 is
   component MultTable_Freq300_uid2147 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2148_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2147
      port map ( X => Xtable_c21,
                 Y => Y1_copy2148_c21);
   Y1_c21 <= Y1_copy2148_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2150
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2150 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2150 is
   component MultTable_Freq300_uid2152 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2153_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2152
      port map ( X => Xtable_c21,
                 Y => Y1_copy2153_c21);
   Y1_c21 <= Y1_copy2153_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2155
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2155 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2155 is
   component MultTable_Freq300_uid2157 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2158_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2157
      port map ( X => Xtable_c21,
                 Y => Y1_copy2158_c21);
   Y1_c21 <= Y1_copy2158_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--             IntMultiplierLUT_4_signedx1_signed_Freq300_uid2160
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4_signedx1_signed_Freq300_uid2160 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4_signedx1_signed_Freq300_uid2160 is
   component MultTable_Freq300_uid2162 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2163_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2162
      port map ( X => Xtable_c21,
                 Y => Y1_copy2163_c21);
   Y1_c21 <= Y1_copy2163_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid2165
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid2165 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid2165 is
   component MultTable_Freq300_uid2167 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2168_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2167
      port map ( X => Xtable_c21,
                 Y => Y1_copy2168_c21);
   Y1_c21 <= Y1_copy2168_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_4x1_signed_Freq300_uid2170
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid2170 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid2170 is
   component MultTable_Freq300_uid2172 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2173_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2172
      port map ( X => Xtable_c21,
                 Y => Y1_copy2173_c21);
   Y1_c21 <= Y1_copy2173_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_3_signedx2_Freq300_uid2175
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid2175 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid2175 is
   component MultTable_Freq300_uid2177 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2178_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2177
      port map ( X => Xtable_c21,
                 Y => Y1_copy2178_c21);
   Y1_c21 <= Y1_copy2178_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2180
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2180 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2180 is
   component MultTable_Freq300_uid2182 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2183_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2182
      port map ( X => Xtable_c21,
                 Y => Y1_copy2183_c21);
   Y1_c21 <= Y1_copy2183_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2185
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2185 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2185 is
   component MultTable_Freq300_uid2187 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2188_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2187
      port map ( X => Xtable_c21,
                 Y => Y1_copy2188_c21);
   Y1_c21 <= Y1_copy2188_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2190
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2190 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2190 is
   component MultTable_Freq300_uid2192 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2193_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2192
      port map ( X => Xtable_c21,
                 Y => Y1_copy2193_c21);
   Y1_c21 <= Y1_copy2193_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_3_signedx2_Freq300_uid2195
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid2195 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid2195 is
   component MultTable_Freq300_uid2197 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2198_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2197
      port map ( X => Xtable_c21,
                 Y => Y1_copy2198_c21);
   Y1_c21 <= Y1_copy2198_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2200
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2200 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2200 is
   component MultTable_Freq300_uid2202 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2203_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2202
      port map ( X => Xtable_c21,
                 Y => Y1_copy2203_c21);
   Y1_c21 <= Y1_copy2203_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2205
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2205 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2205 is
   component MultTable_Freq300_uid2207 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2208_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2207
      port map ( X => Xtable_c21,
                 Y => Y1_copy2208_c21);
   Y1_c21 <= Y1_copy2208_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2210
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2210 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2210 is
   component MultTable_Freq300_uid2212 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2213_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2212
      port map ( X => Xtable_c21,
                 Y => Y1_copy2213_c21);
   Y1_c21 <= Y1_copy2213_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_3_signedx2_Freq300_uid2215
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid2215 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid2215 is
   component MultTable_Freq300_uid2217 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2218_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2217
      port map ( X => Xtable_c21,
                 Y => Y1_copy2218_c21);
   Y1_c21 <= Y1_copy2218_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2220
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2220 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2220 is
   component MultTable_Freq300_uid2222 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2223_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2222
      port map ( X => Xtable_c21,
                 Y => Y1_copy2223_c21);
   Y1_c21 <= Y1_copy2223_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2225
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2225 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2225 is
   component MultTable_Freq300_uid2227 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2228_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2227
      port map ( X => Xtable_c21,
                 Y => Y1_copy2228_c21);
   Y1_c21 <= Y1_copy2228_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2230
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2230 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2230 is
   component MultTable_Freq300_uid2232 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2233_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2232
      port map ( X => Xtable_c21,
                 Y => Y1_copy2233_c21);
   Y1_c21 <= Y1_copy2233_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplierLUT_3_signedx2_Freq300_uid2235
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid2235 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid2235 is
   component MultTable_Freq300_uid2237 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2238_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2237
      port map ( X => Xtable_c21,
                 Y => Y1_copy2238_c21);
   Y1_c21 <= Y1_copy2238_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2240
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2240 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2240 is
   component MultTable_Freq300_uid2242 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2243_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2242
      port map ( X => Xtable_c21,
                 Y => Y1_copy2243_c21);
   Y1_c21 <= Y1_copy2243_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2245
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2245 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2245 is
   component MultTable_Freq300_uid2247 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2248_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2247
      port map ( X => Xtable_c21,
                 Y => Y1_copy2248_c21);
   Y1_c21 <= Y1_copy2248_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2250
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2250 is
    port (clk, ce_20, ce_21 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2250 is
   component MultTable_Freq300_uid2252 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c21 :  std_logic_vector(4 downto 0);
signal Y1_c21 :  std_logic_vector(4 downto 0);
signal Y1_copy2253_c21 :  std_logic_vector(4 downto 0);
signal X_c20, X_c21 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               X_c20 <= X;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
            end if;
         end if;
      end process;
Xtable_c21 <= Y & X_c21;
   R <= Y1_c21;
   TableMult: MultTable_Freq300_uid2252
      port map ( X => Xtable_c21,
                 Y => Y1_copy2253_c21);
   Y1_c21 <= Y1_copy2253_c21; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_45_Freq300_uid2580
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_45_Freq300_uid2580 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          X : in  std_logic_vector(44 downto 0);
          Y : in  std_logic_vector(44 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(44 downto 0)   );
end entity;

architecture arch of IntAdder_45_Freq300_uid2580 is
signal Rtmp_c23 :  std_logic_vector(44 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19, Cin_c20, Cin_c21, Cin_c22, Cin_c23 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               Cin_c19 <= Cin_c18;
            end if;
            if ce_20 = '1' then
               Cin_c20 <= Cin_c19;
            end if;
            if ce_21 = '1' then
               Cin_c21 <= Cin_c20;
            end if;
            if ce_22 = '1' then
               Cin_c22 <= Cin_c21;
            end if;
            if ce_23 = '1' then
               Cin_c23 <= Cin_c22;
            end if;
         end if;
      end process;
   Rtmp_c23 <= X + Y + Cin_c23;
   R <= Rtmp_c23;
end architecture;

--------------------------------------------------------------------------------
--    FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid2011
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan, 2012-2014, 2024
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y A
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid2011 is
    port (clk, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          X : in  std_logic_vector(28 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          A : in  std_logic_vector(39 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid2011 is
   component DSPBlock_17x24_Freq300_uid2014 is
      port ( clk, ce_20, ce_21, ce_22 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_12x24_Freq300_uid2016 is
      port ( clk, ce_20, ce_21, ce_22 : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(35 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_signed_Freq300_uid2018 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid2020 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid2025 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid2030 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid2035 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2040 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2045 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2050 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2055 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2060 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2065 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2070 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2075 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2080 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2085 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2090 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2095 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2100 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2105 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2110 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2115 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2120 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2125 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2130 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2135 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2140 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2145 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2150 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2155 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4_signedx1_signed_Freq300_uid2160 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid2165 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid2170 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid2175 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2180 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2185 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2190 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid2195 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2200 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2205 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2210 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid2215 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2220 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2225 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2230 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid2235 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2240 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2245 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2250 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid2256 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid2264 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid2272 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid2288 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid2314 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_45_Freq300_uid2580 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             X : in  std_logic_vector(44 downto 0);
             Y : in  std_logic_vector(44 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(44 downto 0)   );
   end component;

signal XX_c19 :  signed(0+28 downto 0);
signal YY_c21 :  signed(-9+41 downto 0);
signal AA_c19 :  signed(-2+41 downto 0);
signal tile_0_X_c19 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c21 :  std_logic_vector(23 downto 0);
signal tile_0_output_c22 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c22 :  unsigned(40-0 downto 0);
signal bh2012_wm69_0_c22, bh2012_wm69_0_c23 :  std_logic;
signal bh2012_wm68_0_c22, bh2012_wm68_0_c23 :  std_logic;
signal bh2012_wm67_0_c22, bh2012_wm67_0_c23 :  std_logic;
signal bh2012_wm66_0_c22, bh2012_wm66_0_c23 :  std_logic;
signal bh2012_wm65_0_c22, bh2012_wm65_0_c23 :  std_logic;
signal bh2012_wm64_0_c22, bh2012_wm64_0_c23 :  std_logic;
signal bh2012_wm63_0_c22, bh2012_wm63_0_c23 :  std_logic;
signal bh2012_wm62_0_c22, bh2012_wm62_0_c23 :  std_logic;
signal bh2012_wm61_0_c22, bh2012_wm61_0_c23 :  std_logic;
signal bh2012_wm60_0_c22, bh2012_wm60_0_c23 :  std_logic;
signal bh2012_wm59_0_c22, bh2012_wm59_0_c23 :  std_logic;
signal bh2012_wm58_0_c22, bh2012_wm58_0_c23 :  std_logic;
signal bh2012_wm57_0_c22, bh2012_wm57_0_c23 :  std_logic;
signal bh2012_wm56_0_c22, bh2012_wm56_0_c23 :  std_logic;
signal bh2012_wm55_0_c22, bh2012_wm55_0_c23 :  std_logic;
signal bh2012_wm54_0_c22, bh2012_wm54_0_c23 :  std_logic;
signal bh2012_wm53_0_c22, bh2012_wm53_0_c23 :  std_logic;
signal bh2012_wm52_0_c22 :  std_logic;
signal bh2012_wm51_0_c22 :  std_logic;
signal bh2012_wm50_0_c22 :  std_logic;
signal bh2012_wm49_0_c22 :  std_logic;
signal bh2012_wm48_0_c22 :  std_logic;
signal bh2012_wm47_0_c22 :  std_logic;
signal bh2012_wm46_0_c22 :  std_logic;
signal bh2012_wm45_0_c22 :  std_logic;
signal bh2012_wm44_0_c22 :  std_logic;
signal bh2012_wm43_0_c22 :  std_logic;
signal bh2012_wm42_0_c22 :  std_logic;
signal bh2012_wm41_0_c22 :  std_logic;
signal bh2012_wm40_0_c22 :  std_logic;
signal bh2012_wm39_0_c22 :  std_logic;
signal bh2012_wm38_0_c22 :  std_logic;
signal bh2012_wm37_0_c22 :  std_logic;
signal bh2012_wm36_0_c22 :  std_logic;
signal bh2012_wm35_0_c22 :  std_logic;
signal bh2012_wm34_0_c22 :  std_logic;
signal bh2012_wm33_0_c22 :  std_logic;
signal bh2012_wm32_0_c22 :  std_logic;
signal bh2012_wm31_0_c22 :  std_logic;
signal bh2012_wm30_0_c22 :  std_logic;
signal bh2012_wm29_0_c22 :  std_logic;
signal tile_1_X_c19 :  std_logic_vector(11 downto 0);
signal tile_1_Y_c21 :  std_logic_vector(23 downto 0);
signal tile_1_output_c22 :  std_logic_vector(35 downto 0);
signal tile_1_filtered_output_c22 :  signed(35-0 downto 0);
signal bh2012_wm52_1_c22 :  std_logic;
signal bh2012_wm51_1_c22 :  std_logic;
signal bh2012_wm50_1_c22 :  std_logic;
signal bh2012_wm49_1_c22 :  std_logic;
signal bh2012_wm48_1_c22 :  std_logic;
signal bh2012_wm47_1_c22 :  std_logic;
signal bh2012_wm46_1_c22 :  std_logic;
signal bh2012_wm45_1_c22 :  std_logic;
signal bh2012_wm44_1_c22 :  std_logic;
signal bh2012_wm43_1_c22 :  std_logic;
signal bh2012_wm42_1_c22 :  std_logic;
signal bh2012_wm41_1_c22 :  std_logic;
signal bh2012_wm40_1_c22 :  std_logic;
signal bh2012_wm39_1_c22 :  std_logic;
signal bh2012_wm38_1_c22 :  std_logic;
signal bh2012_wm37_1_c22 :  std_logic;
signal bh2012_wm36_1_c22 :  std_logic;
signal bh2012_wm35_1_c22 :  std_logic;
signal bh2012_wm34_1_c22 :  std_logic;
signal bh2012_wm33_1_c22 :  std_logic;
signal bh2012_wm32_1_c22 :  std_logic;
signal bh2012_wm31_1_c22 :  std_logic;
signal bh2012_wm30_1_c22 :  std_logic;
signal bh2012_wm29_1_c22 :  std_logic;
signal bh2012_wm28_0_c22 :  std_logic;
signal bh2012_wm27_0_c22 :  std_logic;
signal bh2012_wm26_0_c22 :  std_logic;
signal bh2012_wm25_0_c22 :  std_logic;
signal bh2012_wm24_0_c22 :  std_logic;
signal bh2012_wm23_0_c22 :  std_logic;
signal bh2012_wm22_0_c22 :  std_logic;
signal bh2012_wm21_0_c22 :  std_logic;
signal bh2012_wm20_0_c22 :  std_logic;
signal bh2012_wm19_0_c22 :  std_logic;
signal bh2012_wm18_0_c22 :  std_logic;
signal bh2012_wm17_0_c22 :  std_logic;
signal tile_2_X_c19 :  std_logic_vector(0 downto 0);
signal tile_2_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_2_output_c21 :  std_logic_vector(0 downto 0);
signal tile_2_filtered_output_c21 :  signed(0-0 downto 0);
signal bh2012_wm21_1_c21, bh2012_wm21_1_c22 :  std_logic;
signal tile_3_X_c19 :  std_logic_vector(3 downto 0);
signal tile_3_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_3_output_c21 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm25_1_c21 :  std_logic;
signal bh2012_wm24_1_c21 :  std_logic;
signal bh2012_wm23_1_c21 :  std_logic;
signal bh2012_wm22_1_c21 :  std_logic;
signal bh2012_wm21_2_c21, bh2012_wm21_2_c22 :  std_logic;
signal tile_4_X_c19 :  std_logic_vector(3 downto 0);
signal tile_4_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_4_output_c21 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm29_2_c21, bh2012_wm29_2_c22 :  std_logic;
signal bh2012_wm28_1_c21, bh2012_wm28_1_c22 :  std_logic;
signal bh2012_wm27_1_c21 :  std_logic;
signal bh2012_wm26_1_c21 :  std_logic;
signal bh2012_wm25_2_c21 :  std_logic;
signal tile_5_X_c19 :  std_logic_vector(3 downto 0);
signal tile_5_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_5_output_c21 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm33_2_c21, bh2012_wm33_2_c22 :  std_logic;
signal bh2012_wm32_2_c21, bh2012_wm32_2_c22 :  std_logic;
signal bh2012_wm31_2_c21, bh2012_wm31_2_c22 :  std_logic;
signal bh2012_wm30_2_c21, bh2012_wm30_2_c22 :  std_logic;
signal bh2012_wm29_3_c21, bh2012_wm29_3_c22 :  std_logic;
signal tile_6_X_c19 :  std_logic_vector(3 downto 0);
signal tile_6_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_6_output_c21 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm37_2_c21, bh2012_wm37_2_c22 :  std_logic;
signal bh2012_wm36_2_c21, bh2012_wm36_2_c22 :  std_logic;
signal bh2012_wm35_2_c21, bh2012_wm35_2_c22 :  std_logic;
signal bh2012_wm34_2_c21, bh2012_wm34_2_c22 :  std_logic;
signal bh2012_wm33_3_c21, bh2012_wm33_3_c22 :  std_logic;
signal tile_7_X_c19 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_7_output_c21 :  std_logic_vector(3 downto 0);
signal tile_7_filtered_output_c21 :  unsigned(3-0 downto 0);
signal bh2012_wm24_2_c21 :  std_logic;
signal bh2012_wm23_2_c21 :  std_logic;
signal bh2012_wm22_2_c21 :  std_logic;
signal bh2012_wm21_3_c21, bh2012_wm21_3_c22 :  std_logic;
signal tile_8_X_c19 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_8_output_c21 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm27_2_c21 :  std_logic;
signal bh2012_wm26_2_c21 :  std_logic;
signal bh2012_wm25_3_c21 :  std_logic;
signal bh2012_wm24_3_c21 :  std_logic;
signal bh2012_wm23_3_c21 :  std_logic;
signal tile_9_X_c19 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_9_output_c21 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm30_3_c21, bh2012_wm30_3_c22 :  std_logic;
signal bh2012_wm29_4_c21, bh2012_wm29_4_c22 :  std_logic;
signal bh2012_wm28_2_c21, bh2012_wm28_2_c22 :  std_logic;
signal bh2012_wm27_3_c21 :  std_logic;
signal bh2012_wm26_3_c21 :  std_logic;
signal tile_10_X_c19 :  std_logic_vector(2 downto 0);
signal tile_10_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_10_output_c21 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm33_4_c21, bh2012_wm33_4_c22 :  std_logic;
signal bh2012_wm32_3_c21, bh2012_wm32_3_c22 :  std_logic;
signal bh2012_wm31_3_c21, bh2012_wm31_3_c22 :  std_logic;
signal bh2012_wm30_4_c21, bh2012_wm30_4_c22 :  std_logic;
signal bh2012_wm29_5_c21, bh2012_wm29_5_c22 :  std_logic;
signal tile_11_X_c19 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_11_output_c21 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm36_3_c21, bh2012_wm36_3_c22 :  std_logic;
signal bh2012_wm35_3_c21, bh2012_wm35_3_c22 :  std_logic;
signal bh2012_wm34_3_c21, bh2012_wm34_3_c22 :  std_logic;
signal bh2012_wm33_5_c21, bh2012_wm33_5_c22 :  std_logic;
signal bh2012_wm32_4_c21, bh2012_wm32_4_c22 :  std_logic;
signal tile_12_X_c19 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_12_output_c21 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm39_2_c21, bh2012_wm39_2_c22 :  std_logic;
signal bh2012_wm38_2_c21 :  std_logic;
signal bh2012_wm37_3_c21, bh2012_wm37_3_c22 :  std_logic;
signal bh2012_wm36_4_c21, bh2012_wm36_4_c22 :  std_logic;
signal bh2012_wm35_4_c21, bh2012_wm35_4_c22 :  std_logic;
signal tile_13_X_c19 :  std_logic_vector(1 downto 0);
signal tile_13_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_13_output_c21 :  std_logic_vector(3 downto 0);
signal tile_13_filtered_output_c21 :  unsigned(3-0 downto 0);
signal bh2012_wm26_4_c21 :  std_logic;
signal bh2012_wm25_4_c21 :  std_logic;
signal bh2012_wm24_4_c21 :  std_logic;
signal bh2012_wm23_4_c21 :  std_logic;
signal tile_14_X_c19 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_14_output_c21 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm29_6_c21 :  std_logic;
signal bh2012_wm28_3_c21, bh2012_wm28_3_c22 :  std_logic;
signal bh2012_wm27_4_c21 :  std_logic;
signal bh2012_wm26_5_c21 :  std_logic;
signal bh2012_wm25_5_c21 :  std_logic;
signal tile_15_X_c19 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_15_output_c21 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm32_5_c21, bh2012_wm32_5_c22 :  std_logic;
signal bh2012_wm31_4_c21, bh2012_wm31_4_c22 :  std_logic;
signal bh2012_wm30_5_c21, bh2012_wm30_5_c22 :  std_logic;
signal bh2012_wm29_7_c21 :  std_logic;
signal bh2012_wm28_4_c21, bh2012_wm28_4_c22 :  std_logic;
signal tile_16_X_c19 :  std_logic_vector(2 downto 0);
signal tile_16_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_16_output_c21 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm35_5_c21, bh2012_wm35_5_c22 :  std_logic;
signal bh2012_wm34_4_c21, bh2012_wm34_4_c22 :  std_logic;
signal bh2012_wm33_6_c21, bh2012_wm33_6_c22 :  std_logic;
signal bh2012_wm32_6_c21 :  std_logic;
signal bh2012_wm31_5_c21, bh2012_wm31_5_c22 :  std_logic;
signal tile_17_X_c19 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_17_output_c21 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm38_3_c21 :  std_logic;
signal bh2012_wm37_4_c21, bh2012_wm37_4_c22 :  std_logic;
signal bh2012_wm36_5_c21, bh2012_wm36_5_c22 :  std_logic;
signal bh2012_wm35_6_c21, bh2012_wm35_6_c22 :  std_logic;
signal bh2012_wm34_5_c21, bh2012_wm34_5_c22 :  std_logic;
signal tile_18_X_c19 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_18_output_c21 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm41_2_c21, bh2012_wm41_2_c22 :  std_logic;
signal bh2012_wm40_2_c21, bh2012_wm40_2_c22 :  std_logic;
signal bh2012_wm39_3_c21, bh2012_wm39_3_c22 :  std_logic;
signal bh2012_wm38_4_c21 :  std_logic;
signal bh2012_wm37_5_c21, bh2012_wm37_5_c22 :  std_logic;
signal tile_19_X_c19 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_19_output_c21 :  std_logic_vector(3 downto 0);
signal tile_19_filtered_output_c21 :  unsigned(3-0 downto 0);
signal bh2012_wm28_5_c21, bh2012_wm28_5_c22 :  std_logic;
signal bh2012_wm27_5_c21 :  std_logic;
signal bh2012_wm26_6_c21 :  std_logic;
signal bh2012_wm25_6_c21 :  std_logic;
signal tile_20_X_c19 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_20_output_c21 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm31_6_c21 :  std_logic;
signal bh2012_wm30_6_c21 :  std_logic;
signal bh2012_wm29_8_c21 :  std_logic;
signal bh2012_wm28_6_c21 :  std_logic;
signal bh2012_wm27_6_c21 :  std_logic;
signal tile_21_X_c19 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_21_output_c21 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm34_6_c21, bh2012_wm34_6_c22 :  std_logic;
signal bh2012_wm33_7_c21, bh2012_wm33_7_c22 :  std_logic;
signal bh2012_wm32_7_c21 :  std_logic;
signal bh2012_wm31_7_c21 :  std_logic;
signal bh2012_wm30_7_c21 :  std_logic;
signal tile_22_X_c19 :  std_logic_vector(2 downto 0);
signal tile_22_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_22_output_c21 :  std_logic_vector(4 downto 0);
signal tile_22_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm37_6_c21 :  std_logic;
signal bh2012_wm36_6_c21, bh2012_wm36_6_c22 :  std_logic;
signal bh2012_wm35_7_c21 :  std_logic;
signal bh2012_wm34_7_c21 :  std_logic;
signal bh2012_wm33_8_c21, bh2012_wm33_8_c22 :  std_logic;
signal tile_23_X_c19 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_23_output_c21 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm40_3_c21, bh2012_wm40_3_c22 :  std_logic;
signal bh2012_wm39_4_c21, bh2012_wm39_4_c22 :  std_logic;
signal bh2012_wm38_5_c21 :  std_logic;
signal bh2012_wm37_7_c21 :  std_logic;
signal bh2012_wm36_7_c21 :  std_logic;
signal tile_24_X_c19 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_24_output_c21 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm43_2_c21, bh2012_wm43_2_c22 :  std_logic;
signal bh2012_wm42_2_c21, bh2012_wm42_2_c22 :  std_logic;
signal bh2012_wm41_3_c21, bh2012_wm41_3_c22 :  std_logic;
signal bh2012_wm40_4_c21, bh2012_wm40_4_c22 :  std_logic;
signal bh2012_wm39_5_c21, bh2012_wm39_5_c22 :  std_logic;
signal tile_25_X_c19 :  std_logic_vector(1 downto 0);
signal tile_25_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_25_output_c21 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c21 :  unsigned(3-0 downto 0);
signal bh2012_wm30_8_c21 :  std_logic;
signal bh2012_wm29_9_c21 :  std_logic;
signal bh2012_wm28_7_c21 :  std_logic;
signal bh2012_wm27_7_c21 :  std_logic;
signal tile_26_X_c19 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_26_output_c21 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm33_9_c21, bh2012_wm33_9_c22 :  std_logic;
signal bh2012_wm32_8_c21 :  std_logic;
signal bh2012_wm31_8_c21 :  std_logic;
signal bh2012_wm30_9_c21 :  std_logic;
signal bh2012_wm29_10_c21 :  std_logic;
signal tile_27_X_c19 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_27_output_c21 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm36_8_c21 :  std_logic;
signal bh2012_wm35_8_c21 :  std_logic;
signal bh2012_wm34_8_c21 :  std_logic;
signal bh2012_wm33_10_c21, bh2012_wm33_10_c22 :  std_logic;
signal bh2012_wm32_9_c21 :  std_logic;
signal tile_28_X_c19 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_28_output_c21 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm39_6_c21 :  std_logic;
signal bh2012_wm38_6_c21 :  std_logic;
signal bh2012_wm37_8_c21 :  std_logic;
signal bh2012_wm36_9_c21 :  std_logic;
signal bh2012_wm35_9_c21 :  std_logic;
signal tile_29_X_c19 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_29_output_c21 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm42_3_c21, bh2012_wm42_3_c22 :  std_logic;
signal bh2012_wm41_4_c21, bh2012_wm41_4_c22 :  std_logic;
signal bh2012_wm40_5_c21, bh2012_wm40_5_c22 :  std_logic;
signal bh2012_wm39_7_c21 :  std_logic;
signal bh2012_wm38_7_c21 :  std_logic;
signal tile_30_X_c19 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_30_output_c21 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm45_2_c21, bh2012_wm45_2_c22 :  std_logic;
signal bh2012_wm44_2_c21, bh2012_wm44_2_c22 :  std_logic;
signal bh2012_wm43_3_c21, bh2012_wm43_3_c22 :  std_logic;
signal bh2012_wm42_4_c21, bh2012_wm42_4_c22 :  std_logic;
signal bh2012_wm41_5_c21, bh2012_wm41_5_c22 :  std_logic;
signal tile_31_X_c19 :  std_logic_vector(3 downto 0);
signal tile_31_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_31_output_c21 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm12_0_c21 :  std_logic;
signal bh2012_wm11_0_c21 :  std_logic;
signal bh2012_wm10_0_c21 :  std_logic;
signal bh2012_wm9_0_c21 :  std_logic;
signal bh2012_wm8_0_c21 :  std_logic;
signal tile_32_X_c19 :  std_logic_vector(3 downto 0);
signal tile_32_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_32_output_c21 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm16_0_c21 :  std_logic;
signal bh2012_wm15_0_c21 :  std_logic;
signal bh2012_wm14_0_c21 :  std_logic;
signal bh2012_wm13_0_c21 :  std_logic;
signal bh2012_wm12_1_c21 :  std_logic;
signal tile_33_X_c19 :  std_logic_vector(3 downto 0);
signal tile_33_Y_c21 :  std_logic_vector(0 downto 0);
signal tile_33_output_c21 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm20_1_c21, bh2012_wm20_1_c22 :  std_logic;
signal bh2012_wm19_1_c21, bh2012_wm19_1_c22 :  std_logic;
signal bh2012_wm18_1_c21 :  std_logic;
signal bh2012_wm17_1_c21, bh2012_wm17_1_c22 :  std_logic;
signal bh2012_wm16_1_c21 :  std_logic;
signal tile_34_X_c19 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_34_output_c21 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm13_1_c21 :  std_logic;
signal bh2012_wm12_2_c21 :  std_logic;
signal bh2012_wm11_1_c21 :  std_logic;
signal bh2012_wm10_1_c21 :  std_logic;
signal bh2012_wm9_1_c21 :  std_logic;
signal tile_35_X_c19 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_35_output_c21 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm16_2_c21 :  std_logic;
signal bh2012_wm15_1_c21 :  std_logic;
signal bh2012_wm14_1_c21 :  std_logic;
signal bh2012_wm13_2_c21 :  std_logic;
signal bh2012_wm12_3_c21 :  std_logic;
signal tile_36_X_c19 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_36_output_c21 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm19_2_c21, bh2012_wm19_2_c22 :  std_logic;
signal bh2012_wm18_2_c21 :  std_logic;
signal bh2012_wm17_2_c21, bh2012_wm17_2_c22 :  std_logic;
signal bh2012_wm16_3_c21 :  std_logic;
signal bh2012_wm15_2_c21 :  std_logic;
signal tile_37_X_c19 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_37_output_c21 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm22_3_c21 :  std_logic;
signal bh2012_wm21_4_c21, bh2012_wm21_4_c22 :  std_logic;
signal bh2012_wm20_2_c21, bh2012_wm20_2_c22 :  std_logic;
signal bh2012_wm19_3_c21, bh2012_wm19_3_c22 :  std_logic;
signal bh2012_wm18_3_c21 :  std_logic;
signal tile_38_X_c19 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_38_output_c21 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm15_3_c21 :  std_logic;
signal bh2012_wm14_2_c21 :  std_logic;
signal bh2012_wm13_3_c21 :  std_logic;
signal bh2012_wm12_4_c21 :  std_logic;
signal bh2012_wm11_2_c21 :  std_logic;
signal tile_39_X_c19 :  std_logic_vector(2 downto 0);
signal tile_39_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_39_output_c21 :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm18_4_c21 :  std_logic;
signal bh2012_wm17_3_c21, bh2012_wm17_3_c22 :  std_logic;
signal bh2012_wm16_4_c21 :  std_logic;
signal bh2012_wm15_4_c21 :  std_logic;
signal bh2012_wm14_3_c21 :  std_logic;
signal tile_40_X_c19 :  std_logic_vector(2 downto 0);
signal tile_40_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_40_output_c21 :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm21_5_c21, bh2012_wm21_5_c22 :  std_logic;
signal bh2012_wm20_3_c21, bh2012_wm20_3_c22 :  std_logic;
signal bh2012_wm19_4_c21, bh2012_wm19_4_c22 :  std_logic;
signal bh2012_wm18_5_c21 :  std_logic;
signal bh2012_wm17_4_c21, bh2012_wm17_4_c22 :  std_logic;
signal tile_41_X_c19 :  std_logic_vector(2 downto 0);
signal tile_41_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_41_output_c21 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm24_5_c21 :  std_logic;
signal bh2012_wm23_5_c21 :  std_logic;
signal bh2012_wm22_4_c21 :  std_logic;
signal bh2012_wm21_6_c21 :  std_logic;
signal bh2012_wm20_4_c21, bh2012_wm20_4_c22 :  std_logic;
signal tile_42_X_c19 :  std_logic_vector(2 downto 0);
signal tile_42_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_42_output_c21 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm17_5_c21, bh2012_wm17_5_c22 :  std_logic;
signal bh2012_wm16_5_c21 :  std_logic;
signal bh2012_wm15_5_c21 :  std_logic;
signal bh2012_wm14_4_c21 :  std_logic;
signal bh2012_wm13_4_c21 :  std_logic;
signal tile_43_X_c19 :  std_logic_vector(2 downto 0);
signal tile_43_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_43_output_c21 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm20_5_c21, bh2012_wm20_5_c22 :  std_logic;
signal bh2012_wm19_5_c21, bh2012_wm19_5_c22 :  std_logic;
signal bh2012_wm18_6_c21 :  std_logic;
signal bh2012_wm17_6_c21 :  std_logic;
signal bh2012_wm16_6_c21 :  std_logic;
signal tile_44_X_c19 :  std_logic_vector(2 downto 0);
signal tile_44_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_44_output_c21 :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm23_6_c21 :  std_logic;
signal bh2012_wm22_5_c21 :  std_logic;
signal bh2012_wm21_7_c21 :  std_logic;
signal bh2012_wm20_6_c21 :  std_logic;
signal bh2012_wm19_6_c21 :  std_logic;
signal tile_45_X_c19 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_45_output_c21 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm26_7_c21 :  std_logic;
signal bh2012_wm25_7_c21 :  std_logic;
signal bh2012_wm24_6_c21 :  std_logic;
signal bh2012_wm23_7_c21 :  std_logic;
signal bh2012_wm22_6_c21 :  std_logic;
signal tile_46_X_c19 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_46_output_c21 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c21 :  signed(4-0 downto 0);
signal bh2012_wm19_7_c21 :  std_logic;
signal bh2012_wm18_7_c21 :  std_logic;
signal bh2012_wm17_7_c21 :  std_logic;
signal bh2012_wm16_7_c21 :  std_logic;
signal bh2012_wm15_6_c21 :  std_logic;
signal tile_47_X_c19 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_47_output_c21 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm22_7_c21 :  std_logic;
signal bh2012_wm21_8_c21 :  std_logic;
signal bh2012_wm20_7_c21 :  std_logic;
signal bh2012_wm19_8_c21 :  std_logic;
signal bh2012_wm18_8_c21 :  std_logic;
signal tile_48_X_c19 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_48_output_c21 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm25_8_c21 :  std_logic;
signal bh2012_wm24_7_c21 :  std_logic;
signal bh2012_wm23_8_c21 :  std_logic;
signal bh2012_wm22_8_c21 :  std_logic;
signal bh2012_wm21_9_c21 :  std_logic;
signal tile_49_X_c19 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c21 :  std_logic_vector(1 downto 0);
signal tile_49_output_c21 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c21 :  unsigned(4-0 downto 0);
signal bh2012_wm28_8_c21 :  std_logic;
signal bh2012_wm27_8_c21 :  std_logic;
signal bh2012_wm26_8_c21 :  std_logic;
signal bh2012_wm25_9_c21 :  std_logic;
signal bh2012_wm24_8_c21 :  std_logic;
signal bh2012_wm41_6_c19, bh2012_wm41_6_c20, bh2012_wm41_6_c21, bh2012_wm41_6_c22 :  std_logic;
signal bh2012_wm40_6_c19, bh2012_wm40_6_c20, bh2012_wm40_6_c21, bh2012_wm40_6_c22 :  std_logic;
signal bh2012_wm39_8_c19, bh2012_wm39_8_c20, bh2012_wm39_8_c21 :  std_logic;
signal bh2012_wm38_8_c19, bh2012_wm38_8_c20, bh2012_wm38_8_c21, bh2012_wm38_8_c22 :  std_logic;
signal bh2012_wm37_9_c19, bh2012_wm37_9_c20, bh2012_wm37_9_c21 :  std_logic;
signal bh2012_wm36_10_c19, bh2012_wm36_10_c20, bh2012_wm36_10_c21 :  std_logic;
signal bh2012_wm35_10_c19, bh2012_wm35_10_c20, bh2012_wm35_10_c21 :  std_logic;
signal bh2012_wm34_9_c19, bh2012_wm34_9_c20, bh2012_wm34_9_c21 :  std_logic;
signal bh2012_wm33_11_c19, bh2012_wm33_11_c20, bh2012_wm33_11_c21, bh2012_wm33_11_c22 :  std_logic;
signal bh2012_wm32_10_c19, bh2012_wm32_10_c20, bh2012_wm32_10_c21 :  std_logic;
signal bh2012_wm31_9_c19, bh2012_wm31_9_c20, bh2012_wm31_9_c21 :  std_logic;
signal bh2012_wm30_10_c19, bh2012_wm30_10_c20, bh2012_wm30_10_c21 :  std_logic;
signal bh2012_wm29_11_c19, bh2012_wm29_11_c20, bh2012_wm29_11_c21 :  std_logic;
signal bh2012_wm28_9_c19, bh2012_wm28_9_c20, bh2012_wm28_9_c21 :  std_logic;
signal bh2012_wm27_9_c19, bh2012_wm27_9_c20, bh2012_wm27_9_c21 :  std_logic;
signal bh2012_wm26_9_c19, bh2012_wm26_9_c20, bh2012_wm26_9_c21 :  std_logic;
signal bh2012_wm25_10_c19, bh2012_wm25_10_c20, bh2012_wm25_10_c21 :  std_logic;
signal bh2012_wm24_9_c19, bh2012_wm24_9_c20, bh2012_wm24_9_c21 :  std_logic;
signal bh2012_wm23_9_c19, bh2012_wm23_9_c20, bh2012_wm23_9_c21 :  std_logic;
signal bh2012_wm22_9_c19, bh2012_wm22_9_c20, bh2012_wm22_9_c21 :  std_logic;
signal bh2012_wm21_10_c19, bh2012_wm21_10_c20, bh2012_wm21_10_c21 :  std_logic;
signal bh2012_wm20_8_c19, bh2012_wm20_8_c20, bh2012_wm20_8_c21 :  std_logic;
signal bh2012_wm19_9_c19, bh2012_wm19_9_c20, bh2012_wm19_9_c21 :  std_logic;
signal bh2012_wm18_9_c19, bh2012_wm18_9_c20, bh2012_wm18_9_c21 :  std_logic;
signal bh2012_wm17_8_c19, bh2012_wm17_8_c20, bh2012_wm17_8_c21 :  std_logic;
signal bh2012_wm16_8_c19, bh2012_wm16_8_c20, bh2012_wm16_8_c21 :  std_logic;
signal bh2012_wm15_7_c19, bh2012_wm15_7_c20, bh2012_wm15_7_c21 :  std_logic;
signal bh2012_wm14_5_c19, bh2012_wm14_5_c20, bh2012_wm14_5_c21 :  std_logic;
signal bh2012_wm13_5_c19, bh2012_wm13_5_c20, bh2012_wm13_5_c21 :  std_logic;
signal bh2012_wm12_5_c19, bh2012_wm12_5_c20, bh2012_wm12_5_c21 :  std_logic;
signal bh2012_wm11_3_c19, bh2012_wm11_3_c20, bh2012_wm11_3_c21 :  std_logic;
signal bh2012_wm10_2_c19, bh2012_wm10_2_c20, bh2012_wm10_2_c21 :  std_logic;
signal bh2012_wm9_2_c19, bh2012_wm9_2_c20, bh2012_wm9_2_c21 :  std_logic;
signal bh2012_wm8_1_c19, bh2012_wm8_1_c20, bh2012_wm8_1_c21 :  std_logic;
signal bh2012_wm7_0_c19 :  std_logic;
signal bh2012_wm6_0_c19 :  std_logic;
signal bh2012_wm5_0_c19 :  std_logic;
signal bh2012_wm4_0_c19 :  std_logic;
signal bh2012_wm3_0_c19 :  std_logic;
signal bh2012_wm2_0_c19 :  std_logic;
signal bh2012_wm42_5_c0, bh2012_wm42_5_c1, bh2012_wm42_5_c2, bh2012_wm42_5_c3, bh2012_wm42_5_c4, bh2012_wm42_5_c5, bh2012_wm42_5_c6, bh2012_wm42_5_c7, bh2012_wm42_5_c8, bh2012_wm42_5_c9, bh2012_wm42_5_c10, bh2012_wm42_5_c11, bh2012_wm42_5_c12, bh2012_wm42_5_c13, bh2012_wm42_5_c14, bh2012_wm42_5_c15, bh2012_wm42_5_c16, bh2012_wm42_5_c17, bh2012_wm42_5_c18, bh2012_wm42_5_c19, bh2012_wm42_5_c20, bh2012_wm42_5_c21, bh2012_wm42_5_c22 :  std_logic;
signal bh2012_wm33_12_c0, bh2012_wm33_12_c1, bh2012_wm33_12_c2, bh2012_wm33_12_c3, bh2012_wm33_12_c4, bh2012_wm33_12_c5, bh2012_wm33_12_c6, bh2012_wm33_12_c7, bh2012_wm33_12_c8, bh2012_wm33_12_c9, bh2012_wm33_12_c10, bh2012_wm33_12_c11, bh2012_wm33_12_c12, bh2012_wm33_12_c13, bh2012_wm33_12_c14, bh2012_wm33_12_c15, bh2012_wm33_12_c16, bh2012_wm33_12_c17, bh2012_wm33_12_c18, bh2012_wm33_12_c19, bh2012_wm33_12_c20, bh2012_wm33_12_c21, bh2012_wm33_12_c22 :  std_logic;
signal bh2012_wm32_11_c0, bh2012_wm32_11_c1, bh2012_wm32_11_c2, bh2012_wm32_11_c3, bh2012_wm32_11_c4, bh2012_wm32_11_c5, bh2012_wm32_11_c6, bh2012_wm32_11_c7, bh2012_wm32_11_c8, bh2012_wm32_11_c9, bh2012_wm32_11_c10, bh2012_wm32_11_c11, bh2012_wm32_11_c12, bh2012_wm32_11_c13, bh2012_wm32_11_c14, bh2012_wm32_11_c15, bh2012_wm32_11_c16, bh2012_wm32_11_c17, bh2012_wm32_11_c18, bh2012_wm32_11_c19, bh2012_wm32_11_c20, bh2012_wm32_11_c21 :  std_logic;
signal bh2012_wm31_10_c0, bh2012_wm31_10_c1, bh2012_wm31_10_c2, bh2012_wm31_10_c3, bh2012_wm31_10_c4, bh2012_wm31_10_c5, bh2012_wm31_10_c6, bh2012_wm31_10_c7, bh2012_wm31_10_c8, bh2012_wm31_10_c9, bh2012_wm31_10_c10, bh2012_wm31_10_c11, bh2012_wm31_10_c12, bh2012_wm31_10_c13, bh2012_wm31_10_c14, bh2012_wm31_10_c15, bh2012_wm31_10_c16, bh2012_wm31_10_c17, bh2012_wm31_10_c18, bh2012_wm31_10_c19, bh2012_wm31_10_c20, bh2012_wm31_10_c21 :  std_logic;
signal bh2012_wm30_11_c0, bh2012_wm30_11_c1, bh2012_wm30_11_c2, bh2012_wm30_11_c3, bh2012_wm30_11_c4, bh2012_wm30_11_c5, bh2012_wm30_11_c6, bh2012_wm30_11_c7, bh2012_wm30_11_c8, bh2012_wm30_11_c9, bh2012_wm30_11_c10, bh2012_wm30_11_c11, bh2012_wm30_11_c12, bh2012_wm30_11_c13, bh2012_wm30_11_c14, bh2012_wm30_11_c15, bh2012_wm30_11_c16, bh2012_wm30_11_c17, bh2012_wm30_11_c18, bh2012_wm30_11_c19, bh2012_wm30_11_c20, bh2012_wm30_11_c21 :  std_logic;
signal bh2012_wm28_10_c0, bh2012_wm28_10_c1, bh2012_wm28_10_c2, bh2012_wm28_10_c3, bh2012_wm28_10_c4, bh2012_wm28_10_c5, bh2012_wm28_10_c6, bh2012_wm28_10_c7, bh2012_wm28_10_c8, bh2012_wm28_10_c9, bh2012_wm28_10_c10, bh2012_wm28_10_c11, bh2012_wm28_10_c12, bh2012_wm28_10_c13, bh2012_wm28_10_c14, bh2012_wm28_10_c15, bh2012_wm28_10_c16, bh2012_wm28_10_c17, bh2012_wm28_10_c18, bh2012_wm28_10_c19, bh2012_wm28_10_c20, bh2012_wm28_10_c21, bh2012_wm28_10_c22 :  std_logic;
signal bh2012_wm27_10_c0, bh2012_wm27_10_c1, bh2012_wm27_10_c2, bh2012_wm27_10_c3, bh2012_wm27_10_c4, bh2012_wm27_10_c5, bh2012_wm27_10_c6, bh2012_wm27_10_c7, bh2012_wm27_10_c8, bh2012_wm27_10_c9, bh2012_wm27_10_c10, bh2012_wm27_10_c11, bh2012_wm27_10_c12, bh2012_wm27_10_c13, bh2012_wm27_10_c14, bh2012_wm27_10_c15, bh2012_wm27_10_c16, bh2012_wm27_10_c17, bh2012_wm27_10_c18, bh2012_wm27_10_c19, bh2012_wm27_10_c20, bh2012_wm27_10_c21 :  std_logic;
signal bh2012_wm26_10_c0, bh2012_wm26_10_c1, bh2012_wm26_10_c2, bh2012_wm26_10_c3, bh2012_wm26_10_c4, bh2012_wm26_10_c5, bh2012_wm26_10_c6, bh2012_wm26_10_c7, bh2012_wm26_10_c8, bh2012_wm26_10_c9, bh2012_wm26_10_c10, bh2012_wm26_10_c11, bh2012_wm26_10_c12, bh2012_wm26_10_c13, bh2012_wm26_10_c14, bh2012_wm26_10_c15, bh2012_wm26_10_c16, bh2012_wm26_10_c17, bh2012_wm26_10_c18, bh2012_wm26_10_c19, bh2012_wm26_10_c20, bh2012_wm26_10_c21 :  std_logic;
signal bh2012_wm24_10_c0, bh2012_wm24_10_c1, bh2012_wm24_10_c2, bh2012_wm24_10_c3, bh2012_wm24_10_c4, bh2012_wm24_10_c5, bh2012_wm24_10_c6, bh2012_wm24_10_c7, bh2012_wm24_10_c8, bh2012_wm24_10_c9, bh2012_wm24_10_c10, bh2012_wm24_10_c11, bh2012_wm24_10_c12, bh2012_wm24_10_c13, bh2012_wm24_10_c14, bh2012_wm24_10_c15, bh2012_wm24_10_c16, bh2012_wm24_10_c17, bh2012_wm24_10_c18, bh2012_wm24_10_c19, bh2012_wm24_10_c20, bh2012_wm24_10_c21 :  std_logic;
signal bh2012_wm23_10_c0, bh2012_wm23_10_c1, bh2012_wm23_10_c2, bh2012_wm23_10_c3, bh2012_wm23_10_c4, bh2012_wm23_10_c5, bh2012_wm23_10_c6, bh2012_wm23_10_c7, bh2012_wm23_10_c8, bh2012_wm23_10_c9, bh2012_wm23_10_c10, bh2012_wm23_10_c11, bh2012_wm23_10_c12, bh2012_wm23_10_c13, bh2012_wm23_10_c14, bh2012_wm23_10_c15, bh2012_wm23_10_c16, bh2012_wm23_10_c17, bh2012_wm23_10_c18, bh2012_wm23_10_c19, bh2012_wm23_10_c20, bh2012_wm23_10_c21 :  std_logic;
signal bh2012_wm22_10_c0, bh2012_wm22_10_c1, bh2012_wm22_10_c2, bh2012_wm22_10_c3, bh2012_wm22_10_c4, bh2012_wm22_10_c5, bh2012_wm22_10_c6, bh2012_wm22_10_c7, bh2012_wm22_10_c8, bh2012_wm22_10_c9, bh2012_wm22_10_c10, bh2012_wm22_10_c11, bh2012_wm22_10_c12, bh2012_wm22_10_c13, bh2012_wm22_10_c14, bh2012_wm22_10_c15, bh2012_wm22_10_c16, bh2012_wm22_10_c17, bh2012_wm22_10_c18, bh2012_wm22_10_c19, bh2012_wm22_10_c20, bh2012_wm22_10_c21, bh2012_wm22_10_c22 :  std_logic;
signal bh2012_wm21_11_c0, bh2012_wm21_11_c1, bh2012_wm21_11_c2, bh2012_wm21_11_c3, bh2012_wm21_11_c4, bh2012_wm21_11_c5, bh2012_wm21_11_c6, bh2012_wm21_11_c7, bh2012_wm21_11_c8, bh2012_wm21_11_c9, bh2012_wm21_11_c10, bh2012_wm21_11_c11, bh2012_wm21_11_c12, bh2012_wm21_11_c13, bh2012_wm21_11_c14, bh2012_wm21_11_c15, bh2012_wm21_11_c16, bh2012_wm21_11_c17, bh2012_wm21_11_c18, bh2012_wm21_11_c19, bh2012_wm21_11_c20, bh2012_wm21_11_c21 :  std_logic;
signal bh2012_wm19_10_c0 :  std_logic;
signal bh2012_wm18_10_c0, bh2012_wm18_10_c1, bh2012_wm18_10_c2, bh2012_wm18_10_c3, bh2012_wm18_10_c4, bh2012_wm18_10_c5, bh2012_wm18_10_c6, bh2012_wm18_10_c7, bh2012_wm18_10_c8, bh2012_wm18_10_c9, bh2012_wm18_10_c10, bh2012_wm18_10_c11, bh2012_wm18_10_c12, bh2012_wm18_10_c13, bh2012_wm18_10_c14, bh2012_wm18_10_c15, bh2012_wm18_10_c16, bh2012_wm18_10_c17, bh2012_wm18_10_c18, bh2012_wm18_10_c19, bh2012_wm18_10_c20, bh2012_wm18_10_c21 :  std_logic;
signal bh2012_wm14_6_c0 :  std_logic;
signal bh2012_wm10_3_c0, bh2012_wm10_3_c1, bh2012_wm10_3_c2, bh2012_wm10_3_c3, bh2012_wm10_3_c4, bh2012_wm10_3_c5, bh2012_wm10_3_c6, bh2012_wm10_3_c7, bh2012_wm10_3_c8, bh2012_wm10_3_c9, bh2012_wm10_3_c10, bh2012_wm10_3_c11, bh2012_wm10_3_c12, bh2012_wm10_3_c13, bh2012_wm10_3_c14, bh2012_wm10_3_c15, bh2012_wm10_3_c16, bh2012_wm10_3_c17, bh2012_wm10_3_c18, bh2012_wm10_3_c19, bh2012_wm10_3_c20, bh2012_wm10_3_c21 :  std_logic;
signal bh2012_wm7_1_c0, bh2012_wm7_1_c1, bh2012_wm7_1_c2, bh2012_wm7_1_c3, bh2012_wm7_1_c4, bh2012_wm7_1_c5, bh2012_wm7_1_c6, bh2012_wm7_1_c7, bh2012_wm7_1_c8, bh2012_wm7_1_c9, bh2012_wm7_1_c10, bh2012_wm7_1_c11, bh2012_wm7_1_c12, bh2012_wm7_1_c13, bh2012_wm7_1_c14, bh2012_wm7_1_c15, bh2012_wm7_1_c16, bh2012_wm7_1_c17, bh2012_wm7_1_c18, bh2012_wm7_1_c19 :  std_logic;
signal bh2012_wm6_1_c0, bh2012_wm6_1_c1, bh2012_wm6_1_c2, bh2012_wm6_1_c3, bh2012_wm6_1_c4, bh2012_wm6_1_c5, bh2012_wm6_1_c6, bh2012_wm6_1_c7, bh2012_wm6_1_c8, bh2012_wm6_1_c9, bh2012_wm6_1_c10, bh2012_wm6_1_c11, bh2012_wm6_1_c12, bh2012_wm6_1_c13, bh2012_wm6_1_c14, bh2012_wm6_1_c15, bh2012_wm6_1_c16, bh2012_wm6_1_c17, bh2012_wm6_1_c18, bh2012_wm6_1_c19 :  std_logic;
signal bh2012_wm5_1_c0, bh2012_wm5_1_c1, bh2012_wm5_1_c2, bh2012_wm5_1_c3, bh2012_wm5_1_c4, bh2012_wm5_1_c5, bh2012_wm5_1_c6, bh2012_wm5_1_c7, bh2012_wm5_1_c8, bh2012_wm5_1_c9, bh2012_wm5_1_c10, bh2012_wm5_1_c11, bh2012_wm5_1_c12, bh2012_wm5_1_c13, bh2012_wm5_1_c14, bh2012_wm5_1_c15, bh2012_wm5_1_c16, bh2012_wm5_1_c17, bh2012_wm5_1_c18, bh2012_wm5_1_c19 :  std_logic;
signal bh2012_wm4_1_c0, bh2012_wm4_1_c1, bh2012_wm4_1_c2, bh2012_wm4_1_c3, bh2012_wm4_1_c4, bh2012_wm4_1_c5, bh2012_wm4_1_c6, bh2012_wm4_1_c7, bh2012_wm4_1_c8, bh2012_wm4_1_c9, bh2012_wm4_1_c10, bh2012_wm4_1_c11, bh2012_wm4_1_c12, bh2012_wm4_1_c13, bh2012_wm4_1_c14, bh2012_wm4_1_c15, bh2012_wm4_1_c16, bh2012_wm4_1_c17, bh2012_wm4_1_c18, bh2012_wm4_1_c19 :  std_logic;
signal bh2012_wm3_1_c0, bh2012_wm3_1_c1, bh2012_wm3_1_c2, bh2012_wm3_1_c3, bh2012_wm3_1_c4, bh2012_wm3_1_c5, bh2012_wm3_1_c6, bh2012_wm3_1_c7, bh2012_wm3_1_c8, bh2012_wm3_1_c9, bh2012_wm3_1_c10, bh2012_wm3_1_c11, bh2012_wm3_1_c12, bh2012_wm3_1_c13, bh2012_wm3_1_c14, bh2012_wm3_1_c15, bh2012_wm3_1_c16, bh2012_wm3_1_c17, bh2012_wm3_1_c18, bh2012_wm3_1_c19 :  std_logic;
signal bh2012_wm1_0_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2257_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2257_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm52_2_c22, bh2012_wm52_2_c23 :  std_logic;
signal bh2012_wm51_2_c22, bh2012_wm51_2_c23 :  std_logic;
signal bh2012_wm50_2_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_copy2258_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2259_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2259_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm50_3_c22 :  std_logic;
signal bh2012_wm49_2_c22 :  std_logic;
signal bh2012_wm48_2_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_copy2260_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2261_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2261_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm48_3_c22 :  std_logic;
signal bh2012_wm47_2_c22 :  std_logic;
signal bh2012_wm46_2_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_copy2262_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2265_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm46_3_c22 :  std_logic;
signal bh2012_wm45_3_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_copy2266_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2267_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2267_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm45_4_c22 :  std_logic;
signal bh2012_wm44_3_c22 :  std_logic;
signal bh2012_wm43_4_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_copy2268_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2269_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm43_5_c22 :  std_logic;
signal bh2012_wm42_6_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_copy2270_c22 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2273_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm42_7_c22 :  std_logic;
signal bh2012_wm41_7_c22 :  std_logic;
signal bh2012_wm40_7_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_copy2274_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2275_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm41_8_c22 :  std_logic;
signal bh2012_wm40_8_c22 :  std_logic;
signal bh2012_wm39_9_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_copy2276_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2277_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm40_9_c22 :  std_logic;
signal bh2012_wm39_10_c22 :  std_logic;
signal bh2012_wm38_9_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_copy2278_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2279_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm39_11_c22 :  std_logic;
signal bh2012_wm38_10_c22 :  std_logic;
signal bh2012_wm37_10_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_copy2280_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In0_c21, Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm39_12_c22 :  std_logic;
signal bh2012_wm38_11_c22 :  std_logic;
signal bh2012_wm37_11_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_copy2282_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2283_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm38_12_c21, bh2012_wm38_12_c22 :  std_logic;
signal bh2012_wm37_12_c21, bh2012_wm37_12_c22 :  std_logic;
signal bh2012_wm36_11_c21 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_copy2284_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2285_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm37_13_c22 :  std_logic;
signal bh2012_wm36_12_c22 :  std_logic;
signal bh2012_wm35_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_copy2286_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm37_14_c22 :  std_logic;
signal bh2012_wm36_13_c22 :  std_logic;
signal bh2012_wm35_12_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_copy2290_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2291_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm36_14_c22 :  std_logic;
signal bh2012_wm35_13_c22 :  std_logic;
signal bh2012_wm34_10_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_copy2292_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm36_15_c22 :  std_logic;
signal bh2012_wm35_14_c22 :  std_logic;
signal bh2012_wm34_11_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_copy2294_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2295_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm35_15_c22 :  std_logic;
signal bh2012_wm34_12_c22 :  std_logic;
signal bh2012_wm33_13_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_copy2296_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm35_16_c22 :  std_logic;
signal bh2012_wm34_13_c22 :  std_logic;
signal bh2012_wm33_14_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_copy2298_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2299_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm34_14_c22 :  std_logic;
signal bh2012_wm33_15_c22 :  std_logic;
signal bh2012_wm32_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_copy2300_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2301_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_c21 :  std_logic_vector(1 downto 0);
signal bh2012_wm34_15_c21, bh2012_wm34_15_c22 :  std_logic;
signal bh2012_wm33_16_c21, bh2012_wm33_16_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_copy2302_c21 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2303_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm33_17_c22 :  std_logic;
signal bh2012_wm32_13_c22 :  std_logic;
signal bh2012_wm31_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_copy2304_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2305_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm33_18_c22 :  std_logic;
signal bh2012_wm32_14_c22 :  std_logic;
signal bh2012_wm31_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_copy2306_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2307_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm32_15_c22 :  std_logic;
signal bh2012_wm31_13_c22 :  std_logic;
signal bh2012_wm30_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_copy2308_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2309_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm32_16_c21, bh2012_wm32_16_c22 :  std_logic;
signal bh2012_wm31_14_c21, bh2012_wm31_14_c22 :  std_logic;
signal bh2012_wm30_13_c21, bh2012_wm30_13_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_copy2310_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2311_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm31_15_c22 :  std_logic;
signal bh2012_wm30_14_c22 :  std_logic;
signal bh2012_wm29_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_copy2312_c22 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2315_In0_c21 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm31_16_c21, bh2012_wm31_16_c22 :  std_logic;
signal bh2012_wm30_15_c21, bh2012_wm30_15_c22 :  std_logic;
signal bh2012_wm29_13_c21, bh2012_wm29_13_c22 :  std_logic;
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_copy2316_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2317_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm30_16_c22 :  std_logic;
signal bh2012_wm29_14_c22 :  std_logic;
signal bh2012_wm28_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_copy2318_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2319_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm30_17_c21, bh2012_wm30_17_c22 :  std_logic;
signal bh2012_wm29_15_c21, bh2012_wm29_15_c22 :  std_logic;
signal bh2012_wm28_12_c21, bh2012_wm28_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_copy2320_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2321_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm29_16_c22 :  std_logic;
signal bh2012_wm28_13_c22 :  std_logic;
signal bh2012_wm27_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_copy2322_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2323_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm29_17_c21, bh2012_wm29_17_c22 :  std_logic;
signal bh2012_wm28_14_c21, bh2012_wm28_14_c22 :  std_logic;
signal bh2012_wm27_12_c21, bh2012_wm27_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_copy2324_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2325_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm28_15_c22 :  std_logic;
signal bh2012_wm27_13_c22 :  std_logic;
signal bh2012_wm26_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_copy2326_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm28_16_c22 :  std_logic;
signal bh2012_wm27_14_c22 :  std_logic;
signal bh2012_wm26_12_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_copy2328_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2329_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm27_15_c21, bh2012_wm27_15_c22 :  std_logic;
signal bh2012_wm26_13_c21, bh2012_wm26_13_c22 :  std_logic;
signal bh2012_wm25_11_c21, bh2012_wm25_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_copy2330_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm27_16_c22 :  std_logic;
signal bh2012_wm26_14_c22 :  std_logic;
signal bh2012_wm25_12_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_copy2332_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2333_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm26_15_c21, bh2012_wm26_15_c22 :  std_logic;
signal bh2012_wm25_13_c21, bh2012_wm25_13_c22 :  std_logic;
signal bh2012_wm24_11_c21, bh2012_wm24_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_copy2334_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm26_16_c22 :  std_logic;
signal bh2012_wm25_14_c22 :  std_logic;
signal bh2012_wm24_12_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_copy2336_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2337_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm25_15_c21, bh2012_wm25_15_c22 :  std_logic;
signal bh2012_wm24_13_c21, bh2012_wm24_13_c22 :  std_logic;
signal bh2012_wm23_11_c21, bh2012_wm23_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_copy2338_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm25_16_c22 :  std_logic;
signal bh2012_wm24_14_c22 :  std_logic;
signal bh2012_wm23_12_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_copy2340_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2341_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm24_15_c21, bh2012_wm24_15_c22 :  std_logic;
signal bh2012_wm23_13_c21, bh2012_wm23_13_c22 :  std_logic;
signal bh2012_wm22_11_c21, bh2012_wm22_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_copy2342_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm24_16_c22 :  std_logic;
signal bh2012_wm23_14_c22 :  std_logic;
signal bh2012_wm22_12_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_copy2344_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2345_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm23_15_c21, bh2012_wm23_15_c22 :  std_logic;
signal bh2012_wm22_13_c21, bh2012_wm22_13_c22 :  std_logic;
signal bh2012_wm21_12_c21, bh2012_wm21_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_copy2346_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm23_16_c22 :  std_logic;
signal bh2012_wm22_14_c22 :  std_logic;
signal bh2012_wm21_13_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_copy2348_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2349_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm22_15_c21, bh2012_wm22_15_c22 :  std_logic;
signal bh2012_wm21_14_c21, bh2012_wm21_14_c22 :  std_logic;
signal bh2012_wm20_9_c21, bh2012_wm20_9_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_copy2350_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2351_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_c21 :  std_logic_vector(1 downto 0);
signal bh2012_wm22_16_c21, bh2012_wm22_16_c22 :  std_logic;
signal bh2012_wm21_15_c21, bh2012_wm21_15_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_copy2352_c21 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2353_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm21_16_c22 :  std_logic;
signal bh2012_wm20_10_c22 :  std_logic;
signal bh2012_wm19_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_copy2354_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2355_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm21_17_c21, bh2012_wm21_17_c22 :  std_logic;
signal bh2012_wm20_11_c21, bh2012_wm20_11_c22 :  std_logic;
signal bh2012_wm19_12_c21, bh2012_wm19_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_copy2356_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2357_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm20_12_c22 :  std_logic;
signal bh2012_wm19_13_c22 :  std_logic;
signal bh2012_wm18_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_copy2358_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2359_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_c21 :  std_logic_vector(1 downto 0);
signal bh2012_wm20_13_c21, bh2012_wm20_13_c22 :  std_logic;
signal bh2012_wm19_14_c21, bh2012_wm19_14_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_copy2360_c21 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2361_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm19_15_c22 :  std_logic;
signal bh2012_wm18_12_c22 :  std_logic;
signal bh2012_wm17_9_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_copy2362_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In0_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm19_16_c22 :  std_logic;
signal bh2012_wm18_13_c22 :  std_logic;
signal bh2012_wm17_10_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_copy2364_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2365_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm18_14_c21, bh2012_wm18_14_c22 :  std_logic;
signal bh2012_wm17_11_c21, bh2012_wm17_11_c22 :  std_logic;
signal bh2012_wm16_9_c21, bh2012_wm16_9_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_copy2366_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In0_c21 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c21 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm18_15_c21, bh2012_wm18_15_c22 :  std_logic;
signal bh2012_wm17_12_c21, bh2012_wm17_12_c22 :  std_logic;
signal bh2012_wm16_10_c21, bh2012_wm16_10_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_copy2368_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2369_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm17_13_c22 :  std_logic;
signal bh2012_wm16_11_c22 :  std_logic;
signal bh2012_wm15_8_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_copy2370_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2371_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_c21 :  std_logic_vector(1 downto 0);
signal bh2012_wm17_14_c21, bh2012_wm17_14_c22 :  std_logic;
signal bh2012_wm16_12_c21, bh2012_wm16_12_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_copy2372_c21 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2373_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm16_13_c21, bh2012_wm16_13_c22 :  std_logic;
signal bh2012_wm15_9_c21, bh2012_wm15_9_c22 :  std_logic;
signal bh2012_wm14_7_c21 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_copy2374_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2375_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2375_In1_c21 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm16_14_c21, bh2012_wm16_14_c22 :  std_logic;
signal bh2012_wm15_10_c21, bh2012_wm15_10_c22 :  std_logic;
signal bh2012_wm14_8_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_copy2376_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2377_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm15_11_c21, bh2012_wm15_11_c22 :  std_logic;
signal bh2012_wm14_9_c21 :  std_logic;
signal bh2012_wm13_6_c21 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_copy2378_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2379_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm14_10_c21 :  std_logic;
signal bh2012_wm13_7_c21 :  std_logic;
signal bh2012_wm12_6_c21 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_copy2380_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2381_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm13_8_c21 :  std_logic;
signal bh2012_wm12_7_c21 :  std_logic;
signal bh2012_wm11_4_c21 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_copy2382_c21 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2383_In0_c21 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm12_8_c21 :  std_logic;
signal bh2012_wm11_5_c21 :  std_logic;
signal bh2012_wm10_4_c21 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_copy2384_c21 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2385_In0_c21 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2385_In1_c21 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm11_6_c21, bh2012_wm11_6_c22 :  std_logic;
signal bh2012_wm10_5_c21 :  std_logic;
signal bh2012_wm9_3_c21 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_copy2386_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2387_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2387_In1_c21 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm10_6_c21 :  std_logic;
signal bh2012_wm9_4_c21, bh2012_wm9_4_c22 :  std_logic;
signal bh2012_wm8_2_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_copy2388_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c19, Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c20, Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c21 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_c21 :  std_logic_vector(2 downto 0);
signal bh2012_wm8_3_c21 :  std_logic;
signal bh2012_wm7_2_c21 :  std_logic;
signal bh2012_wm6_2_c21 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_copy2390_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2391_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2391_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh2012_wm6_3_c19, bh2012_wm6_3_c20, bh2012_wm6_3_c21 :  std_logic;
signal bh2012_wm5_2_c19 :  std_logic;
signal bh2012_wm4_2_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_copy2392_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2393_In0_c19 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2393_In1_c19 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh2012_wm4_3_c19 :  std_logic;
signal bh2012_wm3_2_c19 :  std_logic;
signal bh2012_wm2_1_c19 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_copy2394_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2395_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2395_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm50_4_c22, bh2012_wm50_4_c23 :  std_logic;
signal bh2012_wm49_3_c22, bh2012_wm49_3_c23 :  std_logic;
signal bh2012_wm48_4_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_copy2396_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2397_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2397_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm48_5_c22 :  std_logic;
signal bh2012_wm47_3_c22 :  std_logic;
signal bh2012_wm46_4_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_copy2398_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2399_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2399_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm46_5_c22 :  std_logic;
signal bh2012_wm45_5_c22 :  std_logic;
signal bh2012_wm44_4_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_copy2400_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2401_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm44_5_c22 :  std_logic;
signal bh2012_wm43_6_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_copy2402_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2403_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2403_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm43_7_c22 :  std_logic;
signal bh2012_wm42_8_c22 :  std_logic;
signal bh2012_wm41_9_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_copy2404_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2405_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm41_10_c22 :  std_logic;
signal bh2012_wm40_10_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_copy2406_c22 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2407_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2407_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm40_11_c22 :  std_logic;
signal bh2012_wm39_13_c22 :  std_logic;
signal bh2012_wm38_13_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_copy2408_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2409_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm39_14_c22 :  std_logic;
signal bh2012_wm38_14_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_copy2410_c22 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2411_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2411_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm38_15_c22 :  std_logic;
signal bh2012_wm37_15_c22 :  std_logic;
signal bh2012_wm36_16_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_copy2412_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm37_16_c22 :  std_logic;
signal bh2012_wm36_17_c22 :  std_logic;
signal bh2012_wm35_17_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_copy2414_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2415_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm36_18_c22 :  std_logic;
signal bh2012_wm35_18_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_copy2416_c22 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2417_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm35_19_c22 :  std_logic;
signal bh2012_wm34_16_c22 :  std_logic;
signal bh2012_wm33_19_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_copy2418_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2419_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm34_17_c22 :  std_logic;
signal bh2012_wm33_20_c22 :  std_logic;
signal bh2012_wm32_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_copy2420_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2421_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm33_21_c22 :  std_logic;
signal bh2012_wm32_18_c22 :  std_logic;
signal bh2012_wm31_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_copy2422_c22 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2423_In0_c22 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm32_19_c22 :  std_logic;
signal bh2012_wm31_18_c22 :  std_logic;
signal bh2012_wm30_18_c22 :  std_logic;
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_copy2424_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2425_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm31_19_c22 :  std_logic;
signal bh2012_wm30_19_c22 :  std_logic;
signal bh2012_wm29_18_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_copy2426_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2427_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm30_20_c22, bh2012_wm30_20_c23 :  std_logic;
signal bh2012_wm29_19_c22 :  std_logic;
signal bh2012_wm28_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_copy2428_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2429_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm29_20_c22 :  std_logic;
signal bh2012_wm28_18_c22 :  std_logic;
signal bh2012_wm27_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_copy2430_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2431_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm28_19_c22 :  std_logic;
signal bh2012_wm27_18_c22 :  std_logic;
signal bh2012_wm26_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_copy2432_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2433_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm27_19_c22 :  std_logic;
signal bh2012_wm26_18_c22 :  std_logic;
signal bh2012_wm25_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_copy2434_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2435_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm26_19_c22 :  std_logic;
signal bh2012_wm25_18_c22 :  std_logic;
signal bh2012_wm24_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_copy2436_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2437_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm25_19_c22, bh2012_wm25_19_c23 :  std_logic;
signal bh2012_wm24_18_c22 :  std_logic;
signal bh2012_wm23_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_copy2438_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2439_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm24_19_c22 :  std_logic;
signal bh2012_wm23_18_c22 :  std_logic;
signal bh2012_wm22_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_copy2440_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2441_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm23_19_c22, bh2012_wm23_19_c23 :  std_logic;
signal bh2012_wm22_18_c22 :  std_logic;
signal bh2012_wm21_18_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_copy2442_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2443_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm22_19_c22 :  std_logic;
signal bh2012_wm21_19_c22 :  std_logic;
signal bh2012_wm20_14_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_copy2444_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2445_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm21_20_c22 :  std_logic;
signal bh2012_wm20_15_c22 :  std_logic;
signal bh2012_wm19_17_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_copy2446_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm20_16_c22 :  std_logic;
signal bh2012_wm19_18_c22 :  std_logic;
signal bh2012_wm18_16_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_copy2448_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2449_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm19_19_c22 :  std_logic;
signal bh2012_wm18_17_c22 :  std_logic;
signal bh2012_wm17_15_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_copy2450_c22 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2451_In0_c22 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm18_18_c22 :  std_logic;
signal bh2012_wm17_16_c22 :  std_logic;
signal bh2012_wm16_15_c22 :  std_logic;
signal Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_copy2452_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2453_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm17_17_c22, bh2012_wm17_17_c23 :  std_logic;
signal bh2012_wm16_16_c22 :  std_logic;
signal bh2012_wm15_12_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_copy2454_c22 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2455_In0_c22 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm16_17_c22 :  std_logic;
signal bh2012_wm15_13_c22 :  std_logic;
signal bh2012_wm14_11_c22 :  std_logic;
signal Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_copy2456_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm15_14_c22, bh2012_wm15_14_c23 :  std_logic;
signal bh2012_wm14_12_c22 :  std_logic;
signal bh2012_wm13_9_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_copy2458_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In0_c21 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c21 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm14_13_c22 :  std_logic;
signal bh2012_wm13_10_c22 :  std_logic;
signal bh2012_wm12_9_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_copy2460_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_copy2460_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2461_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm13_11_c22, bh2012_wm13_11_c23 :  std_logic;
signal bh2012_wm12_10_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_copy2462_c21, Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_copy2462_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2463_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2463_In1_c21 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm12_11_c22 :  std_logic;
signal bh2012_wm11_7_c22 :  std_logic;
signal bh2012_wm10_7_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_copy2464_c21, Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_copy2464_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2465_In0_c21 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2465_In1_c21 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm10_8_c22 :  std_logic;
signal bh2012_wm9_5_c22 :  std_logic;
signal bh2012_wm8_4_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_copy2466_c21, Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_copy2466_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2467_In0_c21 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2467_In1_c21 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm8_5_c22 :  std_logic;
signal bh2012_wm7_3_c22 :  std_logic;
signal bh2012_wm6_4_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_copy2468_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_copy2468_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In0_c21 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c21 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm6_5_c22 :  std_logic;
signal bh2012_wm5_3_c22 :  std_logic;
signal bh2012_wm4_4_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_copy2470_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_copy2470_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2471_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2471_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh2012_wm4_5_c19, bh2012_wm4_5_c20, bh2012_wm4_5_c21, bh2012_wm4_5_c22 :  std_logic;
signal bh2012_wm3_3_c19 :  std_logic;
signal bh2012_wm2_2_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_copy2472_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh2012_wm2_3_c19 :  std_logic;
signal bh2012_wm1_1_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_copy2474_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2475_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2475_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm48_6_c22, bh2012_wm48_6_c23 :  std_logic;
signal bh2012_wm47_4_c22, bh2012_wm47_4_c23 :  std_logic;
signal bh2012_wm46_6_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_copy2476_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2477_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2477_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm46_7_c22 :  std_logic;
signal bh2012_wm45_6_c22 :  std_logic;
signal bh2012_wm44_6_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_copy2478_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2479_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2479_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm44_7_c22 :  std_logic;
signal bh2012_wm43_8_c22 :  std_logic;
signal bh2012_wm42_9_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_copy2480_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2481_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2481_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm41_11_c22 :  std_logic;
signal bh2012_wm40_12_c22, bh2012_wm40_12_c23 :  std_logic;
signal bh2012_wm39_15_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_copy2482_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2483_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_c22 :  std_logic_vector(1 downto 0);
signal bh2012_wm39_16_c22 :  std_logic;
signal bh2012_wm38_16_c22 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_copy2484_c22 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2485_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2485_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm38_17_c22 :  std_logic;
signal bh2012_wm37_17_c22 :  std_logic;
signal bh2012_wm36_19_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_copy2486_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm36_20_c22 :  std_logic;
signal bh2012_wm35_20_c22, bh2012_wm35_20_c23 :  std_logic;
signal bh2012_wm34_18_c22, bh2012_wm34_18_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_copy2488_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2489_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2489_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm35_21_c23 :  std_logic;
signal bh2012_wm34_19_c23 :  std_logic;
signal bh2012_wm33_22_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_copy2490_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_copy2490_c23 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm33_23_c23 :  std_logic;
signal bh2012_wm32_20_c23 :  std_logic;
signal bh2012_wm31_20_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_copy2492_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_copy2492_c23 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2493_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_c23 :  std_logic_vector(1 downto 0);
signal bh2012_wm32_21_c23 :  std_logic;
signal bh2012_wm31_21_c23 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_copy2494_c22, Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_copy2494_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2495_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2495_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm31_22_c23 :  std_logic;
signal bh2012_wm30_21_c23 :  std_logic;
signal bh2012_wm29_21_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_copy2496_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_copy2496_c23 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2497_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_c23 :  std_logic_vector(1 downto 0);
signal bh2012_wm29_22_c23 :  std_logic;
signal bh2012_wm28_20_c23 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_copy2498_c22, Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_copy2498_c23 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm28_21_c23 :  std_logic;
signal bh2012_wm27_20_c23 :  std_logic;
signal bh2012_wm26_20_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_copy2500_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_copy2500_c23 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2501_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_c23 :  std_logic_vector(1 downto 0);
signal bh2012_wm27_21_c23 :  std_logic;
signal bh2012_wm26_21_c23 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_copy2502_c22, Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_copy2502_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2503_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2503_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm26_22_c23 :  std_logic;
signal bh2012_wm25_20_c23 :  std_logic;
signal bh2012_wm24_20_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_copy2504_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_copy2504_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2505_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2505_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm24_21_c23 :  std_logic;
signal bh2012_wm23_20_c23 :  std_logic;
signal bh2012_wm22_20_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_copy2506_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_copy2506_c23 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm22_21_c22, bh2012_wm22_21_c23 :  std_logic;
signal bh2012_wm21_21_c22, bh2012_wm21_21_c23 :  std_logic;
signal bh2012_wm20_17_c22, bh2012_wm20_17_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_copy2508_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2509_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_c23 :  std_logic_vector(1 downto 0);
signal bh2012_wm21_22_c23 :  std_logic;
signal bh2012_wm20_18_c23 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_copy2510_c22, Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_copy2510_c23 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c0, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c1, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c2, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c3, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c4, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c5, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c6, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c7, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c8, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c9, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c10, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c11, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c12, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c13, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c14, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c15, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c16, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c17, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c18, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm20_19_c23 :  std_logic;
signal bh2012_wm19_20_c23 :  std_logic;
signal bh2012_wm18_19_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_copy2512_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_copy2512_c23 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2513_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_c23 :  std_logic_vector(1 downto 0);
signal bh2012_wm19_21_c23 :  std_logic;
signal bh2012_wm18_20_c23 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_copy2514_c22, Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_copy2514_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2515_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2515_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm18_21_c23 :  std_logic;
signal bh2012_wm17_18_c23 :  std_logic;
signal bh2012_wm16_18_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_copy2516_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_copy2516_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2517_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2517_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm16_19_c23 :  std_logic;
signal bh2012_wm15_15_c23 :  std_logic;
signal bh2012_wm14_14_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_copy2518_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_copy2518_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2519_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2519_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm14_15_c23 :  std_logic;
signal bh2012_wm13_12_c23 :  std_logic;
signal bh2012_wm12_12_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_copy2520_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_copy2520_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2521_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2521_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm12_13_c22, bh2012_wm12_13_c23 :  std_logic;
signal bh2012_wm11_8_c22 :  std_logic;
signal bh2012_wm10_9_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_copy2522_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2523_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2523_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm10_10_c22 :  std_logic;
signal bh2012_wm9_6_c22 :  std_logic;
signal bh2012_wm8_6_c22 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_copy2524_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2525_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2525_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm8_7_c22 :  std_logic;
signal bh2012_wm7_4_c22 :  std_logic;
signal bh2012_wm6_6_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_copy2526_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2527_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2527_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm6_7_c22 :  std_logic;
signal bh2012_wm5_4_c22 :  std_logic;
signal bh2012_wm4_6_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_copy2528_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm4_7_c22 :  std_logic;
signal bh2012_wm3_4_c22 :  std_logic;
signal bh2012_wm2_4_c22 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_copy2530_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2531_In0_c19 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2531_In1_c19 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_c19 :  std_logic_vector(2 downto 0);
signal bh2012_wm2_5_c19, bh2012_wm2_5_c20, bh2012_wm2_5_c21, bh2012_wm2_5_c22 :  std_logic;
signal bh2012_wm1_2_c19 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_copy2532_c19 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2533_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2533_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm46_8_c23 :  std_logic;
signal bh2012_wm45_7_c23 :  std_logic;
signal bh2012_wm44_8_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_copy2534_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_copy2534_c23 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2535_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2535_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm44_9_c23 :  std_logic;
signal bh2012_wm43_9_c23 :  std_logic;
signal bh2012_wm42_10_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_copy2536_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_copy2536_c23 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2537_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2537_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm42_11_c23 :  std_logic;
signal bh2012_wm41_12_c23 :  std_logic;
signal bh2012_wm40_13_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_copy2538_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_copy2538_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2539_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2539_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm39_17_c23 :  std_logic;
signal bh2012_wm38_18_c23 :  std_logic;
signal bh2012_wm37_18_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_copy2540_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_copy2540_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2541_In0_c22 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2541_In1_c22 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm37_19_c23 :  std_logic;
signal bh2012_wm36_21_c23 :  std_logic;
signal bh2012_wm35_22_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_copy2542_c22, Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_copy2542_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2543_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2543_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm35_23_c23 :  std_logic;
signal bh2012_wm34_20_c23 :  std_logic;
signal bh2012_wm33_24_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_copy2544_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2545_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2545_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm33_25_c23 :  std_logic;
signal bh2012_wm32_22_c23 :  std_logic;
signal bh2012_wm31_23_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_copy2546_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2547_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2547_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm31_24_c23 :  std_logic;
signal bh2012_wm30_22_c23 :  std_logic;
signal bh2012_wm29_23_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_copy2548_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2549_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2549_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm29_24_c23 :  std_logic;
signal bh2012_wm28_22_c23 :  std_logic;
signal bh2012_wm27_22_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_copy2550_c23 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2551_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_c23 :  std_logic_vector(1 downto 0);
signal bh2012_wm27_23_c23 :  std_logic;
signal bh2012_wm26_23_c23 :  std_logic;
signal Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_copy2552_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2553_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2553_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm26_24_c23 :  std_logic;
signal bh2012_wm25_21_c23 :  std_logic;
signal bh2012_wm24_22_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_copy2554_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2555_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2555_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm24_23_c23 :  std_logic;
signal bh2012_wm23_21_c23 :  std_logic;
signal bh2012_wm22_22_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_copy2556_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2557_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2557_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm22_23_c23 :  std_logic;
signal bh2012_wm21_23_c23 :  std_logic;
signal bh2012_wm20_20_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_copy2558_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2559_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2559_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm20_21_c23 :  std_logic;
signal bh2012_wm19_22_c23 :  std_logic;
signal bh2012_wm18_22_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_copy2560_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2561_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2561_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm18_23_c23 :  std_logic;
signal bh2012_wm17_19_c23 :  std_logic;
signal bh2012_wm16_20_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_copy2562_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2563_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2563_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm16_21_c23 :  std_logic;
signal bh2012_wm15_16_c23 :  std_logic;
signal bh2012_wm14_16_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_copy2564_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2565_In0_c23 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2565_In1_c23 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm14_17_c23 :  std_logic;
signal bh2012_wm13_13_c23 :  std_logic;
signal bh2012_wm12_14_c23 :  std_logic;
signal Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_copy2566_c23 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In0_c23 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In1_c22, Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In1_c23 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_c23 :  std_logic_vector(2 downto 0);
signal bh2012_wm12_15_c23 :  std_logic;
signal bh2012_wm11_9_c23 :  std_logic;
signal bh2012_wm10_11_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_copy2568_c23 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2569_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2569_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm10_12_c22, bh2012_wm10_12_c23 :  std_logic;
signal bh2012_wm9_7_c22, bh2012_wm9_7_c23 :  std_logic;
signal bh2012_wm8_8_c22, bh2012_wm8_8_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_copy2570_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2571_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2571_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm8_9_c22, bh2012_wm8_9_c23 :  std_logic;
signal bh2012_wm7_5_c22, bh2012_wm7_5_c23 :  std_logic;
signal bh2012_wm6_8_c22, bh2012_wm6_8_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_copy2572_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2573_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2573_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm6_9_c22, bh2012_wm6_9_c23 :  std_logic;
signal bh2012_wm5_5_c22, bh2012_wm5_5_c23 :  std_logic;
signal bh2012_wm4_8_c22, bh2012_wm4_8_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_copy2574_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2575_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2575_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm4_9_c22, bh2012_wm4_9_c23 :  std_logic;
signal bh2012_wm3_5_c22, bh2012_wm3_5_c23 :  std_logic;
signal bh2012_wm2_6_c22, bh2012_wm2_6_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_copy2576_c22 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In0_c22 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c19, Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c20, Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c21, Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c22 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_c22 :  std_logic_vector(2 downto 0);
signal bh2012_wm2_7_c22, bh2012_wm2_7_c23 :  std_logic;
signal bh2012_wm1_3_c22, bh2012_wm1_3_c23 :  std_logic;
signal Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_copy2578_c22 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh2012_24_c23 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh2012_In0_c23 :  std_logic_vector(44 downto 0);
signal bitheapFinalAdd_bh2012_In1_c23 :  std_logic_vector(44 downto 0);
signal bitheapFinalAdd_bh2012_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh2012_Out_c23 :  std_logic_vector(44 downto 0);
signal bitheapResult_bh2012_c23 :  std_logic_vector(68 downto 0);
signal RR_c23 :  signed(-1+41 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
               bh2012_wm41_6_c20 <= bh2012_wm41_6_c19;
               bh2012_wm40_6_c20 <= bh2012_wm40_6_c19;
               bh2012_wm39_8_c20 <= bh2012_wm39_8_c19;
               bh2012_wm38_8_c20 <= bh2012_wm38_8_c19;
               bh2012_wm37_9_c20 <= bh2012_wm37_9_c19;
               bh2012_wm36_10_c20 <= bh2012_wm36_10_c19;
               bh2012_wm35_10_c20 <= bh2012_wm35_10_c19;
               bh2012_wm34_9_c20 <= bh2012_wm34_9_c19;
               bh2012_wm33_11_c20 <= bh2012_wm33_11_c19;
               bh2012_wm32_10_c20 <= bh2012_wm32_10_c19;
               bh2012_wm31_9_c20 <= bh2012_wm31_9_c19;
               bh2012_wm30_10_c20 <= bh2012_wm30_10_c19;
               bh2012_wm29_11_c20 <= bh2012_wm29_11_c19;
               bh2012_wm28_9_c20 <= bh2012_wm28_9_c19;
               bh2012_wm27_9_c20 <= bh2012_wm27_9_c19;
               bh2012_wm26_9_c20 <= bh2012_wm26_9_c19;
               bh2012_wm25_10_c20 <= bh2012_wm25_10_c19;
               bh2012_wm24_9_c20 <= bh2012_wm24_9_c19;
               bh2012_wm23_9_c20 <= bh2012_wm23_9_c19;
               bh2012_wm22_9_c20 <= bh2012_wm22_9_c19;
               bh2012_wm21_10_c20 <= bh2012_wm21_10_c19;
               bh2012_wm20_8_c20 <= bh2012_wm20_8_c19;
               bh2012_wm19_9_c20 <= bh2012_wm19_9_c19;
               bh2012_wm18_9_c20 <= bh2012_wm18_9_c19;
               bh2012_wm17_8_c20 <= bh2012_wm17_8_c19;
               bh2012_wm16_8_c20 <= bh2012_wm16_8_c19;
               bh2012_wm15_7_c20 <= bh2012_wm15_7_c19;
               bh2012_wm14_5_c20 <= bh2012_wm14_5_c19;
               bh2012_wm13_5_c20 <= bh2012_wm13_5_c19;
               bh2012_wm12_5_c20 <= bh2012_wm12_5_c19;
               bh2012_wm11_3_c20 <= bh2012_wm11_3_c19;
               bh2012_wm10_2_c20 <= bh2012_wm10_2_c19;
               bh2012_wm9_2_c20 <= bh2012_wm9_2_c19;
               bh2012_wm8_1_c20 <= bh2012_wm8_1_c19;
               bh2012_wm42_5_c20 <= bh2012_wm42_5_c19;
               bh2012_wm33_12_c20 <= bh2012_wm33_12_c19;
               bh2012_wm32_11_c20 <= bh2012_wm32_11_c19;
               bh2012_wm31_10_c20 <= bh2012_wm31_10_c19;
               bh2012_wm30_11_c20 <= bh2012_wm30_11_c19;
               bh2012_wm28_10_c20 <= bh2012_wm28_10_c19;
               bh2012_wm27_10_c20 <= bh2012_wm27_10_c19;
               bh2012_wm26_10_c20 <= bh2012_wm26_10_c19;
               bh2012_wm24_10_c20 <= bh2012_wm24_10_c19;
               bh2012_wm23_10_c20 <= bh2012_wm23_10_c19;
               bh2012_wm22_10_c20 <= bh2012_wm22_10_c19;
               bh2012_wm21_11_c20 <= bh2012_wm21_11_c19;
               bh2012_wm18_10_c20 <= bh2012_wm18_10_c19;
               bh2012_wm10_3_c20 <= bh2012_wm10_3_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c19;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c20 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c19;
               bh2012_wm6_3_c20 <= bh2012_wm6_3_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c19;
               bh2012_wm4_5_c20 <= bh2012_wm4_5_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c19;
               bh2012_wm2_5_c20 <= bh2012_wm2_5_c19;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c20 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c19;
            end if;
            if ce_21 = '1' then
               bh2012_wm41_6_c21 <= bh2012_wm41_6_c20;
               bh2012_wm40_6_c21 <= bh2012_wm40_6_c20;
               bh2012_wm39_8_c21 <= bh2012_wm39_8_c20;
               bh2012_wm38_8_c21 <= bh2012_wm38_8_c20;
               bh2012_wm37_9_c21 <= bh2012_wm37_9_c20;
               bh2012_wm36_10_c21 <= bh2012_wm36_10_c20;
               bh2012_wm35_10_c21 <= bh2012_wm35_10_c20;
               bh2012_wm34_9_c21 <= bh2012_wm34_9_c20;
               bh2012_wm33_11_c21 <= bh2012_wm33_11_c20;
               bh2012_wm32_10_c21 <= bh2012_wm32_10_c20;
               bh2012_wm31_9_c21 <= bh2012_wm31_9_c20;
               bh2012_wm30_10_c21 <= bh2012_wm30_10_c20;
               bh2012_wm29_11_c21 <= bh2012_wm29_11_c20;
               bh2012_wm28_9_c21 <= bh2012_wm28_9_c20;
               bh2012_wm27_9_c21 <= bh2012_wm27_9_c20;
               bh2012_wm26_9_c21 <= bh2012_wm26_9_c20;
               bh2012_wm25_10_c21 <= bh2012_wm25_10_c20;
               bh2012_wm24_9_c21 <= bh2012_wm24_9_c20;
               bh2012_wm23_9_c21 <= bh2012_wm23_9_c20;
               bh2012_wm22_9_c21 <= bh2012_wm22_9_c20;
               bh2012_wm21_10_c21 <= bh2012_wm21_10_c20;
               bh2012_wm20_8_c21 <= bh2012_wm20_8_c20;
               bh2012_wm19_9_c21 <= bh2012_wm19_9_c20;
               bh2012_wm18_9_c21 <= bh2012_wm18_9_c20;
               bh2012_wm17_8_c21 <= bh2012_wm17_8_c20;
               bh2012_wm16_8_c21 <= bh2012_wm16_8_c20;
               bh2012_wm15_7_c21 <= bh2012_wm15_7_c20;
               bh2012_wm14_5_c21 <= bh2012_wm14_5_c20;
               bh2012_wm13_5_c21 <= bh2012_wm13_5_c20;
               bh2012_wm12_5_c21 <= bh2012_wm12_5_c20;
               bh2012_wm11_3_c21 <= bh2012_wm11_3_c20;
               bh2012_wm10_2_c21 <= bh2012_wm10_2_c20;
               bh2012_wm9_2_c21 <= bh2012_wm9_2_c20;
               bh2012_wm8_1_c21 <= bh2012_wm8_1_c20;
               bh2012_wm42_5_c21 <= bh2012_wm42_5_c20;
               bh2012_wm33_12_c21 <= bh2012_wm33_12_c20;
               bh2012_wm32_11_c21 <= bh2012_wm32_11_c20;
               bh2012_wm31_10_c21 <= bh2012_wm31_10_c20;
               bh2012_wm30_11_c21 <= bh2012_wm30_11_c20;
               bh2012_wm28_10_c21 <= bh2012_wm28_10_c20;
               bh2012_wm27_10_c21 <= bh2012_wm27_10_c20;
               bh2012_wm26_10_c21 <= bh2012_wm26_10_c20;
               bh2012_wm24_10_c21 <= bh2012_wm24_10_c20;
               bh2012_wm23_10_c21 <= bh2012_wm23_10_c20;
               bh2012_wm22_10_c21 <= bh2012_wm22_10_c20;
               bh2012_wm21_11_c21 <= bh2012_wm21_11_c20;
               bh2012_wm18_10_c21 <= bh2012_wm18_10_c20;
               bh2012_wm10_3_c21 <= bh2012_wm10_3_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c20;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c20;
               bh2012_wm6_3_c21 <= bh2012_wm6_3_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c20;
               bh2012_wm4_5_c21 <= bh2012_wm4_5_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c20;
               bh2012_wm2_5_c21 <= bh2012_wm2_5_c20;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c20;
            end if;
            if ce_22 = '1' then
               bh2012_wm21_1_c22 <= bh2012_wm21_1_c21;
               bh2012_wm21_2_c22 <= bh2012_wm21_2_c21;
               bh2012_wm29_2_c22 <= bh2012_wm29_2_c21;
               bh2012_wm28_1_c22 <= bh2012_wm28_1_c21;
               bh2012_wm33_2_c22 <= bh2012_wm33_2_c21;
               bh2012_wm32_2_c22 <= bh2012_wm32_2_c21;
               bh2012_wm31_2_c22 <= bh2012_wm31_2_c21;
               bh2012_wm30_2_c22 <= bh2012_wm30_2_c21;
               bh2012_wm29_3_c22 <= bh2012_wm29_3_c21;
               bh2012_wm37_2_c22 <= bh2012_wm37_2_c21;
               bh2012_wm36_2_c22 <= bh2012_wm36_2_c21;
               bh2012_wm35_2_c22 <= bh2012_wm35_2_c21;
               bh2012_wm34_2_c22 <= bh2012_wm34_2_c21;
               bh2012_wm33_3_c22 <= bh2012_wm33_3_c21;
               bh2012_wm21_3_c22 <= bh2012_wm21_3_c21;
               bh2012_wm30_3_c22 <= bh2012_wm30_3_c21;
               bh2012_wm29_4_c22 <= bh2012_wm29_4_c21;
               bh2012_wm28_2_c22 <= bh2012_wm28_2_c21;
               bh2012_wm33_4_c22 <= bh2012_wm33_4_c21;
               bh2012_wm32_3_c22 <= bh2012_wm32_3_c21;
               bh2012_wm31_3_c22 <= bh2012_wm31_3_c21;
               bh2012_wm30_4_c22 <= bh2012_wm30_4_c21;
               bh2012_wm29_5_c22 <= bh2012_wm29_5_c21;
               bh2012_wm36_3_c22 <= bh2012_wm36_3_c21;
               bh2012_wm35_3_c22 <= bh2012_wm35_3_c21;
               bh2012_wm34_3_c22 <= bh2012_wm34_3_c21;
               bh2012_wm33_5_c22 <= bh2012_wm33_5_c21;
               bh2012_wm32_4_c22 <= bh2012_wm32_4_c21;
               bh2012_wm39_2_c22 <= bh2012_wm39_2_c21;
               bh2012_wm37_3_c22 <= bh2012_wm37_3_c21;
               bh2012_wm36_4_c22 <= bh2012_wm36_4_c21;
               bh2012_wm35_4_c22 <= bh2012_wm35_4_c21;
               bh2012_wm28_3_c22 <= bh2012_wm28_3_c21;
               bh2012_wm32_5_c22 <= bh2012_wm32_5_c21;
               bh2012_wm31_4_c22 <= bh2012_wm31_4_c21;
               bh2012_wm30_5_c22 <= bh2012_wm30_5_c21;
               bh2012_wm28_4_c22 <= bh2012_wm28_4_c21;
               bh2012_wm35_5_c22 <= bh2012_wm35_5_c21;
               bh2012_wm34_4_c22 <= bh2012_wm34_4_c21;
               bh2012_wm33_6_c22 <= bh2012_wm33_6_c21;
               bh2012_wm31_5_c22 <= bh2012_wm31_5_c21;
               bh2012_wm37_4_c22 <= bh2012_wm37_4_c21;
               bh2012_wm36_5_c22 <= bh2012_wm36_5_c21;
               bh2012_wm35_6_c22 <= bh2012_wm35_6_c21;
               bh2012_wm34_5_c22 <= bh2012_wm34_5_c21;
               bh2012_wm41_2_c22 <= bh2012_wm41_2_c21;
               bh2012_wm40_2_c22 <= bh2012_wm40_2_c21;
               bh2012_wm39_3_c22 <= bh2012_wm39_3_c21;
               bh2012_wm37_5_c22 <= bh2012_wm37_5_c21;
               bh2012_wm28_5_c22 <= bh2012_wm28_5_c21;
               bh2012_wm34_6_c22 <= bh2012_wm34_6_c21;
               bh2012_wm33_7_c22 <= bh2012_wm33_7_c21;
               bh2012_wm36_6_c22 <= bh2012_wm36_6_c21;
               bh2012_wm33_8_c22 <= bh2012_wm33_8_c21;
               bh2012_wm40_3_c22 <= bh2012_wm40_3_c21;
               bh2012_wm39_4_c22 <= bh2012_wm39_4_c21;
               bh2012_wm43_2_c22 <= bh2012_wm43_2_c21;
               bh2012_wm42_2_c22 <= bh2012_wm42_2_c21;
               bh2012_wm41_3_c22 <= bh2012_wm41_3_c21;
               bh2012_wm40_4_c22 <= bh2012_wm40_4_c21;
               bh2012_wm39_5_c22 <= bh2012_wm39_5_c21;
               bh2012_wm33_9_c22 <= bh2012_wm33_9_c21;
               bh2012_wm33_10_c22 <= bh2012_wm33_10_c21;
               bh2012_wm42_3_c22 <= bh2012_wm42_3_c21;
               bh2012_wm41_4_c22 <= bh2012_wm41_4_c21;
               bh2012_wm40_5_c22 <= bh2012_wm40_5_c21;
               bh2012_wm45_2_c22 <= bh2012_wm45_2_c21;
               bh2012_wm44_2_c22 <= bh2012_wm44_2_c21;
               bh2012_wm43_3_c22 <= bh2012_wm43_3_c21;
               bh2012_wm42_4_c22 <= bh2012_wm42_4_c21;
               bh2012_wm41_5_c22 <= bh2012_wm41_5_c21;
               bh2012_wm20_1_c22 <= bh2012_wm20_1_c21;
               bh2012_wm19_1_c22 <= bh2012_wm19_1_c21;
               bh2012_wm17_1_c22 <= bh2012_wm17_1_c21;
               bh2012_wm19_2_c22 <= bh2012_wm19_2_c21;
               bh2012_wm17_2_c22 <= bh2012_wm17_2_c21;
               bh2012_wm21_4_c22 <= bh2012_wm21_4_c21;
               bh2012_wm20_2_c22 <= bh2012_wm20_2_c21;
               bh2012_wm19_3_c22 <= bh2012_wm19_3_c21;
               bh2012_wm17_3_c22 <= bh2012_wm17_3_c21;
               bh2012_wm21_5_c22 <= bh2012_wm21_5_c21;
               bh2012_wm20_3_c22 <= bh2012_wm20_3_c21;
               bh2012_wm19_4_c22 <= bh2012_wm19_4_c21;
               bh2012_wm17_4_c22 <= bh2012_wm17_4_c21;
               bh2012_wm20_4_c22 <= bh2012_wm20_4_c21;
               bh2012_wm17_5_c22 <= bh2012_wm17_5_c21;
               bh2012_wm20_5_c22 <= bh2012_wm20_5_c21;
               bh2012_wm19_5_c22 <= bh2012_wm19_5_c21;
               bh2012_wm41_6_c22 <= bh2012_wm41_6_c21;
               bh2012_wm40_6_c22 <= bh2012_wm40_6_c21;
               bh2012_wm38_8_c22 <= bh2012_wm38_8_c21;
               bh2012_wm33_11_c22 <= bh2012_wm33_11_c21;
               bh2012_wm42_5_c22 <= bh2012_wm42_5_c21;
               bh2012_wm33_12_c22 <= bh2012_wm33_12_c21;
               bh2012_wm28_10_c22 <= bh2012_wm28_10_c21;
               bh2012_wm22_10_c22 <= bh2012_wm22_10_c21;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In0_c21;
               bh2012_wm38_12_c22 <= bh2012_wm38_12_c21;
               bh2012_wm37_12_c22 <= bh2012_wm37_12_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In0_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In0_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In0_c21;
               bh2012_wm34_15_c22 <= bh2012_wm34_15_c21;
               bh2012_wm33_16_c22 <= bh2012_wm33_16_c21;
               bh2012_wm32_16_c22 <= bh2012_wm32_16_c21;
               bh2012_wm31_14_c22 <= bh2012_wm31_14_c21;
               bh2012_wm30_13_c22 <= bh2012_wm30_13_c21;
               bh2012_wm31_16_c22 <= bh2012_wm31_16_c21;
               bh2012_wm30_15_c22 <= bh2012_wm30_15_c21;
               bh2012_wm29_13_c22 <= bh2012_wm29_13_c21;
               bh2012_wm30_17_c22 <= bh2012_wm30_17_c21;
               bh2012_wm29_15_c22 <= bh2012_wm29_15_c21;
               bh2012_wm28_12_c22 <= bh2012_wm28_12_c21;
               bh2012_wm29_17_c22 <= bh2012_wm29_17_c21;
               bh2012_wm28_14_c22 <= bh2012_wm28_14_c21;
               bh2012_wm27_12_c22 <= bh2012_wm27_12_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In0_c21;
               bh2012_wm27_15_c22 <= bh2012_wm27_15_c21;
               bh2012_wm26_13_c22 <= bh2012_wm26_13_c21;
               bh2012_wm25_11_c22 <= bh2012_wm25_11_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In0_c21;
               bh2012_wm26_15_c22 <= bh2012_wm26_15_c21;
               bh2012_wm25_13_c22 <= bh2012_wm25_13_c21;
               bh2012_wm24_11_c22 <= bh2012_wm24_11_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In0_c21;
               bh2012_wm25_15_c22 <= bh2012_wm25_15_c21;
               bh2012_wm24_13_c22 <= bh2012_wm24_13_c21;
               bh2012_wm23_11_c22 <= bh2012_wm23_11_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In0_c21;
               bh2012_wm24_15_c22 <= bh2012_wm24_15_c21;
               bh2012_wm23_13_c22 <= bh2012_wm23_13_c21;
               bh2012_wm22_11_c22 <= bh2012_wm22_11_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In0_c21;
               bh2012_wm23_15_c22 <= bh2012_wm23_15_c21;
               bh2012_wm22_13_c22 <= bh2012_wm22_13_c21;
               bh2012_wm21_12_c22 <= bh2012_wm21_12_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In0_c21;
               bh2012_wm22_15_c22 <= bh2012_wm22_15_c21;
               bh2012_wm21_14_c22 <= bh2012_wm21_14_c21;
               bh2012_wm20_9_c22 <= bh2012_wm20_9_c21;
               bh2012_wm22_16_c22 <= bh2012_wm22_16_c21;
               bh2012_wm21_15_c22 <= bh2012_wm21_15_c21;
               bh2012_wm21_17_c22 <= bh2012_wm21_17_c21;
               bh2012_wm20_11_c22 <= bh2012_wm20_11_c21;
               bh2012_wm19_12_c22 <= bh2012_wm19_12_c21;
               bh2012_wm20_13_c22 <= bh2012_wm20_13_c21;
               bh2012_wm19_14_c22 <= bh2012_wm19_14_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In0_c21;
               bh2012_wm18_14_c22 <= bh2012_wm18_14_c21;
               bh2012_wm17_11_c22 <= bh2012_wm17_11_c21;
               bh2012_wm16_9_c22 <= bh2012_wm16_9_c21;
               bh2012_wm18_15_c22 <= bh2012_wm18_15_c21;
               bh2012_wm17_12_c22 <= bh2012_wm17_12_c21;
               bh2012_wm16_10_c22 <= bh2012_wm16_10_c21;
               bh2012_wm17_14_c22 <= bh2012_wm17_14_c21;
               bh2012_wm16_12_c22 <= bh2012_wm16_12_c21;
               bh2012_wm16_13_c22 <= bh2012_wm16_13_c21;
               bh2012_wm15_9_c22 <= bh2012_wm15_9_c21;
               bh2012_wm16_14_c22 <= bh2012_wm16_14_c21;
               bh2012_wm15_10_c22 <= bh2012_wm15_10_c21;
               bh2012_wm15_11_c22 <= bh2012_wm15_11_c21;
               bh2012_wm11_6_c22 <= bh2012_wm11_6_c21;
               bh2012_wm9_4_c22 <= bh2012_wm9_4_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_copy2460_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_copy2460_c21;
               Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_copy2462_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_copy2462_c21;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_copy2464_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_copy2464_c21;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_copy2466_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_copy2466_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_copy2468_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_copy2468_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_copy2470_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_copy2470_c21;
               bh2012_wm4_5_c22 <= bh2012_wm4_5_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c21;
               bh2012_wm2_5_c22 <= bh2012_wm2_5_c21;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c21;
            end if;
            if ce_23 = '1' then
               bh2012_wm69_0_c23 <= bh2012_wm69_0_c22;
               bh2012_wm68_0_c23 <= bh2012_wm68_0_c22;
               bh2012_wm67_0_c23 <= bh2012_wm67_0_c22;
               bh2012_wm66_0_c23 <= bh2012_wm66_0_c22;
               bh2012_wm65_0_c23 <= bh2012_wm65_0_c22;
               bh2012_wm64_0_c23 <= bh2012_wm64_0_c22;
               bh2012_wm63_0_c23 <= bh2012_wm63_0_c22;
               bh2012_wm62_0_c23 <= bh2012_wm62_0_c22;
               bh2012_wm61_0_c23 <= bh2012_wm61_0_c22;
               bh2012_wm60_0_c23 <= bh2012_wm60_0_c22;
               bh2012_wm59_0_c23 <= bh2012_wm59_0_c22;
               bh2012_wm58_0_c23 <= bh2012_wm58_0_c22;
               bh2012_wm57_0_c23 <= bh2012_wm57_0_c22;
               bh2012_wm56_0_c23 <= bh2012_wm56_0_c22;
               bh2012_wm55_0_c23 <= bh2012_wm55_0_c22;
               bh2012_wm54_0_c23 <= bh2012_wm54_0_c22;
               bh2012_wm53_0_c23 <= bh2012_wm53_0_c22;
               bh2012_wm52_2_c23 <= bh2012_wm52_2_c22;
               bh2012_wm51_2_c23 <= bh2012_wm51_2_c22;
               bh2012_wm50_4_c23 <= bh2012_wm50_4_c22;
               bh2012_wm49_3_c23 <= bh2012_wm49_3_c22;
               bh2012_wm30_20_c23 <= bh2012_wm30_20_c22;
               bh2012_wm25_19_c23 <= bh2012_wm25_19_c22;
               bh2012_wm23_19_c23 <= bh2012_wm23_19_c22;
               bh2012_wm17_17_c23 <= bh2012_wm17_17_c22;
               bh2012_wm15_14_c23 <= bh2012_wm15_14_c22;
               bh2012_wm13_11_c23 <= bh2012_wm13_11_c22;
               bh2012_wm48_6_c23 <= bh2012_wm48_6_c22;
               bh2012_wm47_4_c23 <= bh2012_wm47_4_c22;
               bh2012_wm40_12_c23 <= bh2012_wm40_12_c22;
               bh2012_wm35_20_c23 <= bh2012_wm35_20_c22;
               bh2012_wm34_18_c23 <= bh2012_wm34_18_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_copy2490_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_copy2490_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_copy2492_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_copy2492_c22;
               Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_copy2494_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_copy2494_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_copy2496_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_copy2496_c22;
               Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_copy2498_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_copy2498_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_copy2500_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_copy2500_c22;
               Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_copy2502_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_copy2502_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_copy2504_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_copy2504_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_copy2506_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_copy2506_c22;
               bh2012_wm22_21_c23 <= bh2012_wm22_21_c22;
               bh2012_wm21_21_c23 <= bh2012_wm21_21_c22;
               bh2012_wm20_17_c23 <= bh2012_wm20_17_c22;
               Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_copy2510_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_copy2510_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_copy2512_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_copy2512_c22;
               Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_copy2514_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_copy2514_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_copy2516_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_copy2516_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_copy2518_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_copy2518_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_copy2520_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_copy2520_c22;
               bh2012_wm12_13_c23 <= bh2012_wm12_13_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_copy2534_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_copy2534_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_copy2536_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_copy2536_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_copy2538_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_copy2538_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_copy2540_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_copy2540_c22;
               Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_copy2542_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_copy2542_c22;
               Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In1_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In1_c22;
               bh2012_wm10_12_c23 <= bh2012_wm10_12_c22;
               bh2012_wm9_7_c23 <= bh2012_wm9_7_c22;
               bh2012_wm8_8_c23 <= bh2012_wm8_8_c22;
               bh2012_wm8_9_c23 <= bh2012_wm8_9_c22;
               bh2012_wm7_5_c23 <= bh2012_wm7_5_c22;
               bh2012_wm6_8_c23 <= bh2012_wm6_8_c22;
               bh2012_wm6_9_c23 <= bh2012_wm6_9_c22;
               bh2012_wm5_5_c23 <= bh2012_wm5_5_c22;
               bh2012_wm4_8_c23 <= bh2012_wm4_8_c22;
               bh2012_wm4_9_c23 <= bh2012_wm4_9_c22;
               bh2012_wm3_5_c23 <= bh2012_wm3_5_c22;
               bh2012_wm2_6_c23 <= bh2012_wm2_6_c22;
               bh2012_wm2_7_c23 <= bh2012_wm2_7_c22;
               bh2012_wm1_3_c23 <= bh2012_wm1_3_c22;
            end if;
         end if;
      end process;
XX_c19 <= signed(X);
YY_c21 <= signed(Y);
AA_c19 <= signed(A);
   tile_0_X_c19 <= X(16 downto 0);
   tile_0_Y_c21 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid2014
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 X => tile_0_X_c19,
                 Y => tile_0_Y_c21,
                 R => tile_0_output_c22);

   tile_0_filtered_output_c22 <= unsigned(tile_0_output_c22(40 downto 0));
   bh2012_wm69_0_c22 <= tile_0_filtered_output_c22(0);
   bh2012_wm68_0_c22 <= tile_0_filtered_output_c22(1);
   bh2012_wm67_0_c22 <= tile_0_filtered_output_c22(2);
   bh2012_wm66_0_c22 <= tile_0_filtered_output_c22(3);
   bh2012_wm65_0_c22 <= tile_0_filtered_output_c22(4);
   bh2012_wm64_0_c22 <= tile_0_filtered_output_c22(5);
   bh2012_wm63_0_c22 <= tile_0_filtered_output_c22(6);
   bh2012_wm62_0_c22 <= tile_0_filtered_output_c22(7);
   bh2012_wm61_0_c22 <= tile_0_filtered_output_c22(8);
   bh2012_wm60_0_c22 <= tile_0_filtered_output_c22(9);
   bh2012_wm59_0_c22 <= tile_0_filtered_output_c22(10);
   bh2012_wm58_0_c22 <= tile_0_filtered_output_c22(11);
   bh2012_wm57_0_c22 <= tile_0_filtered_output_c22(12);
   bh2012_wm56_0_c22 <= tile_0_filtered_output_c22(13);
   bh2012_wm55_0_c22 <= tile_0_filtered_output_c22(14);
   bh2012_wm54_0_c22 <= tile_0_filtered_output_c22(15);
   bh2012_wm53_0_c22 <= tile_0_filtered_output_c22(16);
   bh2012_wm52_0_c22 <= tile_0_filtered_output_c22(17);
   bh2012_wm51_0_c22 <= tile_0_filtered_output_c22(18);
   bh2012_wm50_0_c22 <= tile_0_filtered_output_c22(19);
   bh2012_wm49_0_c22 <= tile_0_filtered_output_c22(20);
   bh2012_wm48_0_c22 <= tile_0_filtered_output_c22(21);
   bh2012_wm47_0_c22 <= tile_0_filtered_output_c22(22);
   bh2012_wm46_0_c22 <= tile_0_filtered_output_c22(23);
   bh2012_wm45_0_c22 <= tile_0_filtered_output_c22(24);
   bh2012_wm44_0_c22 <= tile_0_filtered_output_c22(25);
   bh2012_wm43_0_c22 <= tile_0_filtered_output_c22(26);
   bh2012_wm42_0_c22 <= tile_0_filtered_output_c22(27);
   bh2012_wm41_0_c22 <= tile_0_filtered_output_c22(28);
   bh2012_wm40_0_c22 <= tile_0_filtered_output_c22(29);
   bh2012_wm39_0_c22 <= tile_0_filtered_output_c22(30);
   bh2012_wm38_0_c22 <= tile_0_filtered_output_c22(31);
   bh2012_wm37_0_c22 <= tile_0_filtered_output_c22(32);
   bh2012_wm36_0_c22 <= tile_0_filtered_output_c22(33);
   bh2012_wm35_0_c22 <= tile_0_filtered_output_c22(34);
   bh2012_wm34_0_c22 <= tile_0_filtered_output_c22(35);
   bh2012_wm33_0_c22 <= tile_0_filtered_output_c22(36);
   bh2012_wm32_0_c22 <= tile_0_filtered_output_c22(37);
   bh2012_wm31_0_c22 <= tile_0_filtered_output_c22(38);
   bh2012_wm30_0_c22 <= tile_0_filtered_output_c22(39);
   bh2012_wm29_0_c22 <= tile_0_filtered_output_c22(40);
   tile_1_X_c19 <= X(28 downto 17);
   tile_1_Y_c21 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_12x24_Freq300_uid2016
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 X => tile_1_X_c19,
                 Y => tile_1_Y_c21,
                 R => tile_1_output_c22);

   tile_1_filtered_output_c22 <= signed(tile_1_output_c22(35 downto 0));
   bh2012_wm52_1_c22 <= tile_1_filtered_output_c22(0);
   bh2012_wm51_1_c22 <= tile_1_filtered_output_c22(1);
   bh2012_wm50_1_c22 <= tile_1_filtered_output_c22(2);
   bh2012_wm49_1_c22 <= tile_1_filtered_output_c22(3);
   bh2012_wm48_1_c22 <= tile_1_filtered_output_c22(4);
   bh2012_wm47_1_c22 <= tile_1_filtered_output_c22(5);
   bh2012_wm46_1_c22 <= tile_1_filtered_output_c22(6);
   bh2012_wm45_1_c22 <= tile_1_filtered_output_c22(7);
   bh2012_wm44_1_c22 <= tile_1_filtered_output_c22(8);
   bh2012_wm43_1_c22 <= tile_1_filtered_output_c22(9);
   bh2012_wm42_1_c22 <= tile_1_filtered_output_c22(10);
   bh2012_wm41_1_c22 <= tile_1_filtered_output_c22(11);
   bh2012_wm40_1_c22 <= tile_1_filtered_output_c22(12);
   bh2012_wm39_1_c22 <= tile_1_filtered_output_c22(13);
   bh2012_wm38_1_c22 <= tile_1_filtered_output_c22(14);
   bh2012_wm37_1_c22 <= tile_1_filtered_output_c22(15);
   bh2012_wm36_1_c22 <= tile_1_filtered_output_c22(16);
   bh2012_wm35_1_c22 <= tile_1_filtered_output_c22(17);
   bh2012_wm34_1_c22 <= tile_1_filtered_output_c22(18);
   bh2012_wm33_1_c22 <= tile_1_filtered_output_c22(19);
   bh2012_wm32_1_c22 <= tile_1_filtered_output_c22(20);
   bh2012_wm31_1_c22 <= tile_1_filtered_output_c22(21);
   bh2012_wm30_1_c22 <= tile_1_filtered_output_c22(22);
   bh2012_wm29_1_c22 <= tile_1_filtered_output_c22(23);
   bh2012_wm28_0_c22 <= tile_1_filtered_output_c22(24);
   bh2012_wm27_0_c22 <= tile_1_filtered_output_c22(25);
   bh2012_wm26_0_c22 <= tile_1_filtered_output_c22(26);
   bh2012_wm25_0_c22 <= tile_1_filtered_output_c22(27);
   bh2012_wm24_0_c22 <= tile_1_filtered_output_c22(28);
   bh2012_wm23_0_c22 <= tile_1_filtered_output_c22(29);
   bh2012_wm22_0_c22 <= tile_1_filtered_output_c22(30);
   bh2012_wm21_0_c22 <= tile_1_filtered_output_c22(31);
   bh2012_wm20_0_c22 <= tile_1_filtered_output_c22(32);
   bh2012_wm19_0_c22 <= tile_1_filtered_output_c22(33);
   bh2012_wm18_0_c22 <= tile_1_filtered_output_c22(34);
   bh2012_wm17_0_c22 <= not tile_1_filtered_output_c22(35);
   tile_2_X_c19 <= X(16 downto 16);
   tile_2_Y_c21 <= Y(32 downto 32);
   tile_2_mult: IntMultiplierLUT_1x1_signed_Freq300_uid2018
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_2_X_c19,
                 Y => tile_2_Y_c21,
                 R => tile_2_output_c21);

   tile_2_filtered_output_c21 <= signed(tile_2_output_c21(0 downto 0));
   bh2012_wm21_1_c21 <= not tile_2_filtered_output_c21(0);
   tile_3_X_c19 <= X(15 downto 12);
   tile_3_Y_c21 <= Y(32 downto 32);
   tile_3_mult: IntMultiplierLUT_4x1_signed_Freq300_uid2020
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_3_X_c19,
                 Y => tile_3_Y_c21,
                 R => tile_3_output_c21);

   tile_3_filtered_output_c21 <= signed(tile_3_output_c21(4 downto 0));
   bh2012_wm25_1_c21 <= tile_3_filtered_output_c21(0);
   bh2012_wm24_1_c21 <= tile_3_filtered_output_c21(1);
   bh2012_wm23_1_c21 <= tile_3_filtered_output_c21(2);
   bh2012_wm22_1_c21 <= tile_3_filtered_output_c21(3);
   bh2012_wm21_2_c21 <= not tile_3_filtered_output_c21(4);
   tile_4_X_c19 <= X(11 downto 8);
   tile_4_Y_c21 <= Y(32 downto 32);
   tile_4_mult: IntMultiplierLUT_4x1_signed_Freq300_uid2025
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_4_X_c19,
                 Y => tile_4_Y_c21,
                 R => tile_4_output_c21);

   tile_4_filtered_output_c21 <= signed(tile_4_output_c21(4 downto 0));
   bh2012_wm29_2_c21 <= tile_4_filtered_output_c21(0);
   bh2012_wm28_1_c21 <= tile_4_filtered_output_c21(1);
   bh2012_wm27_1_c21 <= tile_4_filtered_output_c21(2);
   bh2012_wm26_1_c21 <= tile_4_filtered_output_c21(3);
   bh2012_wm25_2_c21 <= not tile_4_filtered_output_c21(4);
   tile_5_X_c19 <= X(7 downto 4);
   tile_5_Y_c21 <= Y(32 downto 32);
   tile_5_mult: IntMultiplierLUT_4x1_signed_Freq300_uid2030
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_5_X_c19,
                 Y => tile_5_Y_c21,
                 R => tile_5_output_c21);

   tile_5_filtered_output_c21 <= signed(tile_5_output_c21(4 downto 0));
   bh2012_wm33_2_c21 <= tile_5_filtered_output_c21(0);
   bh2012_wm32_2_c21 <= tile_5_filtered_output_c21(1);
   bh2012_wm31_2_c21 <= tile_5_filtered_output_c21(2);
   bh2012_wm30_2_c21 <= tile_5_filtered_output_c21(3);
   bh2012_wm29_3_c21 <= not tile_5_filtered_output_c21(4);
   tile_6_X_c19 <= X(3 downto 0);
   tile_6_Y_c21 <= Y(32 downto 32);
   tile_6_mult: IntMultiplierLUT_4x1_signed_Freq300_uid2035
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_6_X_c19,
                 Y => tile_6_Y_c21,
                 R => tile_6_output_c21);

   tile_6_filtered_output_c21 <= signed(tile_6_output_c21(4 downto 0));
   bh2012_wm37_2_c21 <= tile_6_filtered_output_c21(0);
   bh2012_wm36_2_c21 <= tile_6_filtered_output_c21(1);
   bh2012_wm35_2_c21 <= tile_6_filtered_output_c21(2);
   bh2012_wm34_2_c21 <= tile_6_filtered_output_c21(3);
   bh2012_wm33_3_c21 <= not tile_6_filtered_output_c21(4);
   tile_7_X_c19 <= X(16 downto 15);
   tile_7_Y_c21 <= Y(31 downto 30);
   tile_7_mult: IntMultiplierLUT_2x2_Freq300_uid2040
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_7_X_c19,
                 Y => tile_7_Y_c21,
                 R => tile_7_output_c21);

   tile_7_filtered_output_c21 <= unsigned(tile_7_output_c21(3 downto 0));
   bh2012_wm24_2_c21 <= tile_7_filtered_output_c21(0);
   bh2012_wm23_2_c21 <= tile_7_filtered_output_c21(1);
   bh2012_wm22_2_c21 <= tile_7_filtered_output_c21(2);
   bh2012_wm21_3_c21 <= tile_7_filtered_output_c21(3);
   tile_8_X_c19 <= X(14 downto 12);
   tile_8_Y_c21 <= Y(31 downto 30);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid2045
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_8_X_c19,
                 Y => tile_8_Y_c21,
                 R => tile_8_output_c21);

   tile_8_filtered_output_c21 <= unsigned(tile_8_output_c21(4 downto 0));
   bh2012_wm27_2_c21 <= tile_8_filtered_output_c21(0);
   bh2012_wm26_2_c21 <= tile_8_filtered_output_c21(1);
   bh2012_wm25_3_c21 <= tile_8_filtered_output_c21(2);
   bh2012_wm24_3_c21 <= tile_8_filtered_output_c21(3);
   bh2012_wm23_3_c21 <= tile_8_filtered_output_c21(4);
   tile_9_X_c19 <= X(11 downto 9);
   tile_9_Y_c21 <= Y(31 downto 30);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid2050
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_9_X_c19,
                 Y => tile_9_Y_c21,
                 R => tile_9_output_c21);

   tile_9_filtered_output_c21 <= unsigned(tile_9_output_c21(4 downto 0));
   bh2012_wm30_3_c21 <= tile_9_filtered_output_c21(0);
   bh2012_wm29_4_c21 <= tile_9_filtered_output_c21(1);
   bh2012_wm28_2_c21 <= tile_9_filtered_output_c21(2);
   bh2012_wm27_3_c21 <= tile_9_filtered_output_c21(3);
   bh2012_wm26_3_c21 <= tile_9_filtered_output_c21(4);
   tile_10_X_c19 <= X(8 downto 6);
   tile_10_Y_c21 <= Y(31 downto 30);
   tile_10_mult: IntMultiplierLUT_3x2_Freq300_uid2055
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_10_X_c19,
                 Y => tile_10_Y_c21,
                 R => tile_10_output_c21);

   tile_10_filtered_output_c21 <= unsigned(tile_10_output_c21(4 downto 0));
   bh2012_wm33_4_c21 <= tile_10_filtered_output_c21(0);
   bh2012_wm32_3_c21 <= tile_10_filtered_output_c21(1);
   bh2012_wm31_3_c21 <= tile_10_filtered_output_c21(2);
   bh2012_wm30_4_c21 <= tile_10_filtered_output_c21(3);
   bh2012_wm29_5_c21 <= tile_10_filtered_output_c21(4);
   tile_11_X_c19 <= X(5 downto 3);
   tile_11_Y_c21 <= Y(31 downto 30);
   tile_11_mult: IntMultiplierLUT_3x2_Freq300_uid2060
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_11_X_c19,
                 Y => tile_11_Y_c21,
                 R => tile_11_output_c21);

   tile_11_filtered_output_c21 <= unsigned(tile_11_output_c21(4 downto 0));
   bh2012_wm36_3_c21 <= tile_11_filtered_output_c21(0);
   bh2012_wm35_3_c21 <= tile_11_filtered_output_c21(1);
   bh2012_wm34_3_c21 <= tile_11_filtered_output_c21(2);
   bh2012_wm33_5_c21 <= tile_11_filtered_output_c21(3);
   bh2012_wm32_4_c21 <= tile_11_filtered_output_c21(4);
   tile_12_X_c19 <= X(2 downto 0);
   tile_12_Y_c21 <= Y(31 downto 30);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid2065
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_12_X_c19,
                 Y => tile_12_Y_c21,
                 R => tile_12_output_c21);

   tile_12_filtered_output_c21 <= unsigned(tile_12_output_c21(4 downto 0));
   bh2012_wm39_2_c21 <= tile_12_filtered_output_c21(0);
   bh2012_wm38_2_c21 <= tile_12_filtered_output_c21(1);
   bh2012_wm37_3_c21 <= tile_12_filtered_output_c21(2);
   bh2012_wm36_4_c21 <= tile_12_filtered_output_c21(3);
   bh2012_wm35_4_c21 <= tile_12_filtered_output_c21(4);
   tile_13_X_c19 <= X(16 downto 15);
   tile_13_Y_c21 <= Y(29 downto 28);
   tile_13_mult: IntMultiplierLUT_2x2_Freq300_uid2070
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_13_X_c19,
                 Y => tile_13_Y_c21,
                 R => tile_13_output_c21);

   tile_13_filtered_output_c21 <= unsigned(tile_13_output_c21(3 downto 0));
   bh2012_wm26_4_c21 <= tile_13_filtered_output_c21(0);
   bh2012_wm25_4_c21 <= tile_13_filtered_output_c21(1);
   bh2012_wm24_4_c21 <= tile_13_filtered_output_c21(2);
   bh2012_wm23_4_c21 <= tile_13_filtered_output_c21(3);
   tile_14_X_c19 <= X(14 downto 12);
   tile_14_Y_c21 <= Y(29 downto 28);
   tile_14_mult: IntMultiplierLUT_3x2_Freq300_uid2075
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_14_X_c19,
                 Y => tile_14_Y_c21,
                 R => tile_14_output_c21);

   tile_14_filtered_output_c21 <= unsigned(tile_14_output_c21(4 downto 0));
   bh2012_wm29_6_c21 <= tile_14_filtered_output_c21(0);
   bh2012_wm28_3_c21 <= tile_14_filtered_output_c21(1);
   bh2012_wm27_4_c21 <= tile_14_filtered_output_c21(2);
   bh2012_wm26_5_c21 <= tile_14_filtered_output_c21(3);
   bh2012_wm25_5_c21 <= tile_14_filtered_output_c21(4);
   tile_15_X_c19 <= X(11 downto 9);
   tile_15_Y_c21 <= Y(29 downto 28);
   tile_15_mult: IntMultiplierLUT_3x2_Freq300_uid2080
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_15_X_c19,
                 Y => tile_15_Y_c21,
                 R => tile_15_output_c21);

   tile_15_filtered_output_c21 <= unsigned(tile_15_output_c21(4 downto 0));
   bh2012_wm32_5_c21 <= tile_15_filtered_output_c21(0);
   bh2012_wm31_4_c21 <= tile_15_filtered_output_c21(1);
   bh2012_wm30_5_c21 <= tile_15_filtered_output_c21(2);
   bh2012_wm29_7_c21 <= tile_15_filtered_output_c21(3);
   bh2012_wm28_4_c21 <= tile_15_filtered_output_c21(4);
   tile_16_X_c19 <= X(8 downto 6);
   tile_16_Y_c21 <= Y(29 downto 28);
   tile_16_mult: IntMultiplierLUT_3x2_Freq300_uid2085
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_16_X_c19,
                 Y => tile_16_Y_c21,
                 R => tile_16_output_c21);

   tile_16_filtered_output_c21 <= unsigned(tile_16_output_c21(4 downto 0));
   bh2012_wm35_5_c21 <= tile_16_filtered_output_c21(0);
   bh2012_wm34_4_c21 <= tile_16_filtered_output_c21(1);
   bh2012_wm33_6_c21 <= tile_16_filtered_output_c21(2);
   bh2012_wm32_6_c21 <= tile_16_filtered_output_c21(3);
   bh2012_wm31_5_c21 <= tile_16_filtered_output_c21(4);
   tile_17_X_c19 <= X(5 downto 3);
   tile_17_Y_c21 <= Y(29 downto 28);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid2090
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_17_X_c19,
                 Y => tile_17_Y_c21,
                 R => tile_17_output_c21);

   tile_17_filtered_output_c21 <= unsigned(tile_17_output_c21(4 downto 0));
   bh2012_wm38_3_c21 <= tile_17_filtered_output_c21(0);
   bh2012_wm37_4_c21 <= tile_17_filtered_output_c21(1);
   bh2012_wm36_5_c21 <= tile_17_filtered_output_c21(2);
   bh2012_wm35_6_c21 <= tile_17_filtered_output_c21(3);
   bh2012_wm34_5_c21 <= tile_17_filtered_output_c21(4);
   tile_18_X_c19 <= X(2 downto 0);
   tile_18_Y_c21 <= Y(29 downto 28);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid2095
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_18_X_c19,
                 Y => tile_18_Y_c21,
                 R => tile_18_output_c21);

   tile_18_filtered_output_c21 <= unsigned(tile_18_output_c21(4 downto 0));
   bh2012_wm41_2_c21 <= tile_18_filtered_output_c21(0);
   bh2012_wm40_2_c21 <= tile_18_filtered_output_c21(1);
   bh2012_wm39_3_c21 <= tile_18_filtered_output_c21(2);
   bh2012_wm38_4_c21 <= tile_18_filtered_output_c21(3);
   bh2012_wm37_5_c21 <= tile_18_filtered_output_c21(4);
   tile_19_X_c19 <= X(16 downto 15);
   tile_19_Y_c21 <= Y(27 downto 26);
   tile_19_mult: IntMultiplierLUT_2x2_Freq300_uid2100
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_19_X_c19,
                 Y => tile_19_Y_c21,
                 R => tile_19_output_c21);

   tile_19_filtered_output_c21 <= unsigned(tile_19_output_c21(3 downto 0));
   bh2012_wm28_5_c21 <= tile_19_filtered_output_c21(0);
   bh2012_wm27_5_c21 <= tile_19_filtered_output_c21(1);
   bh2012_wm26_6_c21 <= tile_19_filtered_output_c21(2);
   bh2012_wm25_6_c21 <= tile_19_filtered_output_c21(3);
   tile_20_X_c19 <= X(14 downto 12);
   tile_20_Y_c21 <= Y(27 downto 26);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid2105
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_20_X_c19,
                 Y => tile_20_Y_c21,
                 R => tile_20_output_c21);

   tile_20_filtered_output_c21 <= unsigned(tile_20_output_c21(4 downto 0));
   bh2012_wm31_6_c21 <= tile_20_filtered_output_c21(0);
   bh2012_wm30_6_c21 <= tile_20_filtered_output_c21(1);
   bh2012_wm29_8_c21 <= tile_20_filtered_output_c21(2);
   bh2012_wm28_6_c21 <= tile_20_filtered_output_c21(3);
   bh2012_wm27_6_c21 <= tile_20_filtered_output_c21(4);
   tile_21_X_c19 <= X(11 downto 9);
   tile_21_Y_c21 <= Y(27 downto 26);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid2110
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_21_X_c19,
                 Y => tile_21_Y_c21,
                 R => tile_21_output_c21);

   tile_21_filtered_output_c21 <= unsigned(tile_21_output_c21(4 downto 0));
   bh2012_wm34_6_c21 <= tile_21_filtered_output_c21(0);
   bh2012_wm33_7_c21 <= tile_21_filtered_output_c21(1);
   bh2012_wm32_7_c21 <= tile_21_filtered_output_c21(2);
   bh2012_wm31_7_c21 <= tile_21_filtered_output_c21(3);
   bh2012_wm30_7_c21 <= tile_21_filtered_output_c21(4);
   tile_22_X_c19 <= X(8 downto 6);
   tile_22_Y_c21 <= Y(27 downto 26);
   tile_22_mult: IntMultiplierLUT_3x2_Freq300_uid2115
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_22_X_c19,
                 Y => tile_22_Y_c21,
                 R => tile_22_output_c21);

   tile_22_filtered_output_c21 <= unsigned(tile_22_output_c21(4 downto 0));
   bh2012_wm37_6_c21 <= tile_22_filtered_output_c21(0);
   bh2012_wm36_6_c21 <= tile_22_filtered_output_c21(1);
   bh2012_wm35_7_c21 <= tile_22_filtered_output_c21(2);
   bh2012_wm34_7_c21 <= tile_22_filtered_output_c21(3);
   bh2012_wm33_8_c21 <= tile_22_filtered_output_c21(4);
   tile_23_X_c19 <= X(5 downto 3);
   tile_23_Y_c21 <= Y(27 downto 26);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid2120
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_23_X_c19,
                 Y => tile_23_Y_c21,
                 R => tile_23_output_c21);

   tile_23_filtered_output_c21 <= unsigned(tile_23_output_c21(4 downto 0));
   bh2012_wm40_3_c21 <= tile_23_filtered_output_c21(0);
   bh2012_wm39_4_c21 <= tile_23_filtered_output_c21(1);
   bh2012_wm38_5_c21 <= tile_23_filtered_output_c21(2);
   bh2012_wm37_7_c21 <= tile_23_filtered_output_c21(3);
   bh2012_wm36_7_c21 <= tile_23_filtered_output_c21(4);
   tile_24_X_c19 <= X(2 downto 0);
   tile_24_Y_c21 <= Y(27 downto 26);
   tile_24_mult: IntMultiplierLUT_3x2_Freq300_uid2125
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_24_X_c19,
                 Y => tile_24_Y_c21,
                 R => tile_24_output_c21);

   tile_24_filtered_output_c21 <= unsigned(tile_24_output_c21(4 downto 0));
   bh2012_wm43_2_c21 <= tile_24_filtered_output_c21(0);
   bh2012_wm42_2_c21 <= tile_24_filtered_output_c21(1);
   bh2012_wm41_3_c21 <= tile_24_filtered_output_c21(2);
   bh2012_wm40_4_c21 <= tile_24_filtered_output_c21(3);
   bh2012_wm39_5_c21 <= tile_24_filtered_output_c21(4);
   tile_25_X_c19 <= X(16 downto 15);
   tile_25_Y_c21 <= Y(25 downto 24);
   tile_25_mult: IntMultiplierLUT_2x2_Freq300_uid2130
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_25_X_c19,
                 Y => tile_25_Y_c21,
                 R => tile_25_output_c21);

   tile_25_filtered_output_c21 <= unsigned(tile_25_output_c21(3 downto 0));
   bh2012_wm30_8_c21 <= tile_25_filtered_output_c21(0);
   bh2012_wm29_9_c21 <= tile_25_filtered_output_c21(1);
   bh2012_wm28_7_c21 <= tile_25_filtered_output_c21(2);
   bh2012_wm27_7_c21 <= tile_25_filtered_output_c21(3);
   tile_26_X_c19 <= X(14 downto 12);
   tile_26_Y_c21 <= Y(25 downto 24);
   tile_26_mult: IntMultiplierLUT_3x2_Freq300_uid2135
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_26_X_c19,
                 Y => tile_26_Y_c21,
                 R => tile_26_output_c21);

   tile_26_filtered_output_c21 <= unsigned(tile_26_output_c21(4 downto 0));
   bh2012_wm33_9_c21 <= tile_26_filtered_output_c21(0);
   bh2012_wm32_8_c21 <= tile_26_filtered_output_c21(1);
   bh2012_wm31_8_c21 <= tile_26_filtered_output_c21(2);
   bh2012_wm30_9_c21 <= tile_26_filtered_output_c21(3);
   bh2012_wm29_10_c21 <= tile_26_filtered_output_c21(4);
   tile_27_X_c19 <= X(11 downto 9);
   tile_27_Y_c21 <= Y(25 downto 24);
   tile_27_mult: IntMultiplierLUT_3x2_Freq300_uid2140
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_27_X_c19,
                 Y => tile_27_Y_c21,
                 R => tile_27_output_c21);

   tile_27_filtered_output_c21 <= unsigned(tile_27_output_c21(4 downto 0));
   bh2012_wm36_8_c21 <= tile_27_filtered_output_c21(0);
   bh2012_wm35_8_c21 <= tile_27_filtered_output_c21(1);
   bh2012_wm34_8_c21 <= tile_27_filtered_output_c21(2);
   bh2012_wm33_10_c21 <= tile_27_filtered_output_c21(3);
   bh2012_wm32_9_c21 <= tile_27_filtered_output_c21(4);
   tile_28_X_c19 <= X(8 downto 6);
   tile_28_Y_c21 <= Y(25 downto 24);
   tile_28_mult: IntMultiplierLUT_3x2_Freq300_uid2145
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_28_X_c19,
                 Y => tile_28_Y_c21,
                 R => tile_28_output_c21);

   tile_28_filtered_output_c21 <= unsigned(tile_28_output_c21(4 downto 0));
   bh2012_wm39_6_c21 <= tile_28_filtered_output_c21(0);
   bh2012_wm38_6_c21 <= tile_28_filtered_output_c21(1);
   bh2012_wm37_8_c21 <= tile_28_filtered_output_c21(2);
   bh2012_wm36_9_c21 <= tile_28_filtered_output_c21(3);
   bh2012_wm35_9_c21 <= tile_28_filtered_output_c21(4);
   tile_29_X_c19 <= X(5 downto 3);
   tile_29_Y_c21 <= Y(25 downto 24);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid2150
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_29_X_c19,
                 Y => tile_29_Y_c21,
                 R => tile_29_output_c21);

   tile_29_filtered_output_c21 <= unsigned(tile_29_output_c21(4 downto 0));
   bh2012_wm42_3_c21 <= tile_29_filtered_output_c21(0);
   bh2012_wm41_4_c21 <= tile_29_filtered_output_c21(1);
   bh2012_wm40_5_c21 <= tile_29_filtered_output_c21(2);
   bh2012_wm39_7_c21 <= tile_29_filtered_output_c21(3);
   bh2012_wm38_7_c21 <= tile_29_filtered_output_c21(4);
   tile_30_X_c19 <= X(2 downto 0);
   tile_30_Y_c21 <= Y(25 downto 24);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid2155
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_30_X_c19,
                 Y => tile_30_Y_c21,
                 R => tile_30_output_c21);

   tile_30_filtered_output_c21 <= unsigned(tile_30_output_c21(4 downto 0));
   bh2012_wm45_2_c21 <= tile_30_filtered_output_c21(0);
   bh2012_wm44_2_c21 <= tile_30_filtered_output_c21(1);
   bh2012_wm43_3_c21 <= tile_30_filtered_output_c21(2);
   bh2012_wm42_4_c21 <= tile_30_filtered_output_c21(3);
   bh2012_wm41_5_c21 <= tile_30_filtered_output_c21(4);
   tile_31_X_c19 <= X(28 downto 25);
   tile_31_Y_c21 <= Y(32 downto 32);
   tile_31_mult: IntMultiplierLUT_4_signedx1_signed_Freq300_uid2160
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_31_X_c19,
                 Y => tile_31_Y_c21,
                 R => tile_31_output_c21);

   tile_31_filtered_output_c21 <= signed(tile_31_output_c21(4 downto 0));
   bh2012_wm12_0_c21 <= tile_31_filtered_output_c21(0);
   bh2012_wm11_0_c21 <= tile_31_filtered_output_c21(1);
   bh2012_wm10_0_c21 <= tile_31_filtered_output_c21(2);
   bh2012_wm9_0_c21 <= tile_31_filtered_output_c21(3);
   bh2012_wm8_0_c21 <= not tile_31_filtered_output_c21(4);
   tile_32_X_c19 <= X(24 downto 21);
   tile_32_Y_c21 <= Y(32 downto 32);
   tile_32_mult: IntMultiplierLUT_4x1_signed_Freq300_uid2165
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_32_X_c19,
                 Y => tile_32_Y_c21,
                 R => tile_32_output_c21);

   tile_32_filtered_output_c21 <= signed(tile_32_output_c21(4 downto 0));
   bh2012_wm16_0_c21 <= tile_32_filtered_output_c21(0);
   bh2012_wm15_0_c21 <= tile_32_filtered_output_c21(1);
   bh2012_wm14_0_c21 <= tile_32_filtered_output_c21(2);
   bh2012_wm13_0_c21 <= tile_32_filtered_output_c21(3);
   bh2012_wm12_1_c21 <= not tile_32_filtered_output_c21(4);
   tile_33_X_c19 <= X(20 downto 17);
   tile_33_Y_c21 <= Y(32 downto 32);
   tile_33_mult: IntMultiplierLUT_4x1_signed_Freq300_uid2170
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_33_X_c19,
                 Y => tile_33_Y_c21,
                 R => tile_33_output_c21);

   tile_33_filtered_output_c21 <= signed(tile_33_output_c21(4 downto 0));
   bh2012_wm20_1_c21 <= tile_33_filtered_output_c21(0);
   bh2012_wm19_1_c21 <= tile_33_filtered_output_c21(1);
   bh2012_wm18_1_c21 <= tile_33_filtered_output_c21(2);
   bh2012_wm17_1_c21 <= tile_33_filtered_output_c21(3);
   bh2012_wm16_1_c21 <= not tile_33_filtered_output_c21(4);
   tile_34_X_c19 <= X(28 downto 26);
   tile_34_Y_c21 <= Y(31 downto 30);
   tile_34_mult: IntMultiplierLUT_3_signedx2_Freq300_uid2175
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_34_X_c19,
                 Y => tile_34_Y_c21,
                 R => tile_34_output_c21);

   tile_34_filtered_output_c21 <= signed(tile_34_output_c21(4 downto 0));
   bh2012_wm13_1_c21 <= tile_34_filtered_output_c21(0);
   bh2012_wm12_2_c21 <= tile_34_filtered_output_c21(1);
   bh2012_wm11_1_c21 <= tile_34_filtered_output_c21(2);
   bh2012_wm10_1_c21 <= tile_34_filtered_output_c21(3);
   bh2012_wm9_1_c21 <= not tile_34_filtered_output_c21(4);
   tile_35_X_c19 <= X(25 downto 23);
   tile_35_Y_c21 <= Y(31 downto 30);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid2180
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_35_X_c19,
                 Y => tile_35_Y_c21,
                 R => tile_35_output_c21);

   tile_35_filtered_output_c21 <= unsigned(tile_35_output_c21(4 downto 0));
   bh2012_wm16_2_c21 <= tile_35_filtered_output_c21(0);
   bh2012_wm15_1_c21 <= tile_35_filtered_output_c21(1);
   bh2012_wm14_1_c21 <= tile_35_filtered_output_c21(2);
   bh2012_wm13_2_c21 <= tile_35_filtered_output_c21(3);
   bh2012_wm12_3_c21 <= tile_35_filtered_output_c21(4);
   tile_36_X_c19 <= X(22 downto 20);
   tile_36_Y_c21 <= Y(31 downto 30);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid2185
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_36_X_c19,
                 Y => tile_36_Y_c21,
                 R => tile_36_output_c21);

   tile_36_filtered_output_c21 <= unsigned(tile_36_output_c21(4 downto 0));
   bh2012_wm19_2_c21 <= tile_36_filtered_output_c21(0);
   bh2012_wm18_2_c21 <= tile_36_filtered_output_c21(1);
   bh2012_wm17_2_c21 <= tile_36_filtered_output_c21(2);
   bh2012_wm16_3_c21 <= tile_36_filtered_output_c21(3);
   bh2012_wm15_2_c21 <= tile_36_filtered_output_c21(4);
   tile_37_X_c19 <= X(19 downto 17);
   tile_37_Y_c21 <= Y(31 downto 30);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid2190
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_37_X_c19,
                 Y => tile_37_Y_c21,
                 R => tile_37_output_c21);

   tile_37_filtered_output_c21 <= unsigned(tile_37_output_c21(4 downto 0));
   bh2012_wm22_3_c21 <= tile_37_filtered_output_c21(0);
   bh2012_wm21_4_c21 <= tile_37_filtered_output_c21(1);
   bh2012_wm20_2_c21 <= tile_37_filtered_output_c21(2);
   bh2012_wm19_3_c21 <= tile_37_filtered_output_c21(3);
   bh2012_wm18_3_c21 <= tile_37_filtered_output_c21(4);
   tile_38_X_c19 <= X(28 downto 26);
   tile_38_Y_c21 <= Y(29 downto 28);
   tile_38_mult: IntMultiplierLUT_3_signedx2_Freq300_uid2195
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_38_X_c19,
                 Y => tile_38_Y_c21,
                 R => tile_38_output_c21);

   tile_38_filtered_output_c21 <= signed(tile_38_output_c21(4 downto 0));
   bh2012_wm15_3_c21 <= tile_38_filtered_output_c21(0);
   bh2012_wm14_2_c21 <= tile_38_filtered_output_c21(1);
   bh2012_wm13_3_c21 <= tile_38_filtered_output_c21(2);
   bh2012_wm12_4_c21 <= tile_38_filtered_output_c21(3);
   bh2012_wm11_2_c21 <= not tile_38_filtered_output_c21(4);
   tile_39_X_c19 <= X(25 downto 23);
   tile_39_Y_c21 <= Y(29 downto 28);
   tile_39_mult: IntMultiplierLUT_3x2_Freq300_uid2200
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_39_X_c19,
                 Y => tile_39_Y_c21,
                 R => tile_39_output_c21);

   tile_39_filtered_output_c21 <= unsigned(tile_39_output_c21(4 downto 0));
   bh2012_wm18_4_c21 <= tile_39_filtered_output_c21(0);
   bh2012_wm17_3_c21 <= tile_39_filtered_output_c21(1);
   bh2012_wm16_4_c21 <= tile_39_filtered_output_c21(2);
   bh2012_wm15_4_c21 <= tile_39_filtered_output_c21(3);
   bh2012_wm14_3_c21 <= tile_39_filtered_output_c21(4);
   tile_40_X_c19 <= X(22 downto 20);
   tile_40_Y_c21 <= Y(29 downto 28);
   tile_40_mult: IntMultiplierLUT_3x2_Freq300_uid2205
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_40_X_c19,
                 Y => tile_40_Y_c21,
                 R => tile_40_output_c21);

   tile_40_filtered_output_c21 <= unsigned(tile_40_output_c21(4 downto 0));
   bh2012_wm21_5_c21 <= tile_40_filtered_output_c21(0);
   bh2012_wm20_3_c21 <= tile_40_filtered_output_c21(1);
   bh2012_wm19_4_c21 <= tile_40_filtered_output_c21(2);
   bh2012_wm18_5_c21 <= tile_40_filtered_output_c21(3);
   bh2012_wm17_4_c21 <= tile_40_filtered_output_c21(4);
   tile_41_X_c19 <= X(19 downto 17);
   tile_41_Y_c21 <= Y(29 downto 28);
   tile_41_mult: IntMultiplierLUT_3x2_Freq300_uid2210
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_41_X_c19,
                 Y => tile_41_Y_c21,
                 R => tile_41_output_c21);

   tile_41_filtered_output_c21 <= unsigned(tile_41_output_c21(4 downto 0));
   bh2012_wm24_5_c21 <= tile_41_filtered_output_c21(0);
   bh2012_wm23_5_c21 <= tile_41_filtered_output_c21(1);
   bh2012_wm22_4_c21 <= tile_41_filtered_output_c21(2);
   bh2012_wm21_6_c21 <= tile_41_filtered_output_c21(3);
   bh2012_wm20_4_c21 <= tile_41_filtered_output_c21(4);
   tile_42_X_c19 <= X(28 downto 26);
   tile_42_Y_c21 <= Y(27 downto 26);
   tile_42_mult: IntMultiplierLUT_3_signedx2_Freq300_uid2215
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_42_X_c19,
                 Y => tile_42_Y_c21,
                 R => tile_42_output_c21);

   tile_42_filtered_output_c21 <= signed(tile_42_output_c21(4 downto 0));
   bh2012_wm17_5_c21 <= tile_42_filtered_output_c21(0);
   bh2012_wm16_5_c21 <= tile_42_filtered_output_c21(1);
   bh2012_wm15_5_c21 <= tile_42_filtered_output_c21(2);
   bh2012_wm14_4_c21 <= tile_42_filtered_output_c21(3);
   bh2012_wm13_4_c21 <= not tile_42_filtered_output_c21(4);
   tile_43_X_c19 <= X(25 downto 23);
   tile_43_Y_c21 <= Y(27 downto 26);
   tile_43_mult: IntMultiplierLUT_3x2_Freq300_uid2220
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_43_X_c19,
                 Y => tile_43_Y_c21,
                 R => tile_43_output_c21);

   tile_43_filtered_output_c21 <= unsigned(tile_43_output_c21(4 downto 0));
   bh2012_wm20_5_c21 <= tile_43_filtered_output_c21(0);
   bh2012_wm19_5_c21 <= tile_43_filtered_output_c21(1);
   bh2012_wm18_6_c21 <= tile_43_filtered_output_c21(2);
   bh2012_wm17_6_c21 <= tile_43_filtered_output_c21(3);
   bh2012_wm16_6_c21 <= tile_43_filtered_output_c21(4);
   tile_44_X_c19 <= X(22 downto 20);
   tile_44_Y_c21 <= Y(27 downto 26);
   tile_44_mult: IntMultiplierLUT_3x2_Freq300_uid2225
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_44_X_c19,
                 Y => tile_44_Y_c21,
                 R => tile_44_output_c21);

   tile_44_filtered_output_c21 <= unsigned(tile_44_output_c21(4 downto 0));
   bh2012_wm23_6_c21 <= tile_44_filtered_output_c21(0);
   bh2012_wm22_5_c21 <= tile_44_filtered_output_c21(1);
   bh2012_wm21_7_c21 <= tile_44_filtered_output_c21(2);
   bh2012_wm20_6_c21 <= tile_44_filtered_output_c21(3);
   bh2012_wm19_6_c21 <= tile_44_filtered_output_c21(4);
   tile_45_X_c19 <= X(19 downto 17);
   tile_45_Y_c21 <= Y(27 downto 26);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid2230
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_45_X_c19,
                 Y => tile_45_Y_c21,
                 R => tile_45_output_c21);

   tile_45_filtered_output_c21 <= unsigned(tile_45_output_c21(4 downto 0));
   bh2012_wm26_7_c21 <= tile_45_filtered_output_c21(0);
   bh2012_wm25_7_c21 <= tile_45_filtered_output_c21(1);
   bh2012_wm24_6_c21 <= tile_45_filtered_output_c21(2);
   bh2012_wm23_7_c21 <= tile_45_filtered_output_c21(3);
   bh2012_wm22_6_c21 <= tile_45_filtered_output_c21(4);
   tile_46_X_c19 <= X(28 downto 26);
   tile_46_Y_c21 <= Y(25 downto 24);
   tile_46_mult: IntMultiplierLUT_3_signedx2_Freq300_uid2235
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_46_X_c19,
                 Y => tile_46_Y_c21,
                 R => tile_46_output_c21);

   tile_46_filtered_output_c21 <= signed(tile_46_output_c21(4 downto 0));
   bh2012_wm19_7_c21 <= tile_46_filtered_output_c21(0);
   bh2012_wm18_7_c21 <= tile_46_filtered_output_c21(1);
   bh2012_wm17_7_c21 <= tile_46_filtered_output_c21(2);
   bh2012_wm16_7_c21 <= tile_46_filtered_output_c21(3);
   bh2012_wm15_6_c21 <= not tile_46_filtered_output_c21(4);
   tile_47_X_c19 <= X(25 downto 23);
   tile_47_Y_c21 <= Y(25 downto 24);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid2240
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_47_X_c19,
                 Y => tile_47_Y_c21,
                 R => tile_47_output_c21);

   tile_47_filtered_output_c21 <= unsigned(tile_47_output_c21(4 downto 0));
   bh2012_wm22_7_c21 <= tile_47_filtered_output_c21(0);
   bh2012_wm21_8_c21 <= tile_47_filtered_output_c21(1);
   bh2012_wm20_7_c21 <= tile_47_filtered_output_c21(2);
   bh2012_wm19_8_c21 <= tile_47_filtered_output_c21(3);
   bh2012_wm18_8_c21 <= tile_47_filtered_output_c21(4);
   tile_48_X_c19 <= X(22 downto 20);
   tile_48_Y_c21 <= Y(25 downto 24);
   tile_48_mult: IntMultiplierLUT_3x2_Freq300_uid2245
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_48_X_c19,
                 Y => tile_48_Y_c21,
                 R => tile_48_output_c21);

   tile_48_filtered_output_c21 <= unsigned(tile_48_output_c21(4 downto 0));
   bh2012_wm25_8_c21 <= tile_48_filtered_output_c21(0);
   bh2012_wm24_7_c21 <= tile_48_filtered_output_c21(1);
   bh2012_wm23_8_c21 <= tile_48_filtered_output_c21(2);
   bh2012_wm22_8_c21 <= tile_48_filtered_output_c21(3);
   bh2012_wm21_9_c21 <= tile_48_filtered_output_c21(4);
   tile_49_X_c19 <= X(19 downto 17);
   tile_49_Y_c21 <= Y(25 downto 24);
   tile_49_mult: IntMultiplierLUT_3x2_Freq300_uid2250
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 X => tile_49_X_c19,
                 Y => tile_49_Y_c21,
                 R => tile_49_output_c21);

   tile_49_filtered_output_c21 <= unsigned(tile_49_output_c21(4 downto 0));
   bh2012_wm28_8_c21 <= tile_49_filtered_output_c21(0);
   bh2012_wm27_8_c21 <= tile_49_filtered_output_c21(1);
   bh2012_wm26_8_c21 <= tile_49_filtered_output_c21(2);
   bh2012_wm25_9_c21 <= tile_49_filtered_output_c21(3);
   bh2012_wm24_8_c21 <= tile_49_filtered_output_c21(4);
   bh2012_wm41_6_c19 <= AA_c19(0);
   bh2012_wm40_6_c19 <= AA_c19(1);
   bh2012_wm39_8_c19 <= AA_c19(2);
   bh2012_wm38_8_c19 <= AA_c19(3);
   bh2012_wm37_9_c19 <= AA_c19(4);
   bh2012_wm36_10_c19 <= AA_c19(5);
   bh2012_wm35_10_c19 <= AA_c19(6);
   bh2012_wm34_9_c19 <= AA_c19(7);
   bh2012_wm33_11_c19 <= AA_c19(8);
   bh2012_wm32_10_c19 <= AA_c19(9);
   bh2012_wm31_9_c19 <= AA_c19(10);
   bh2012_wm30_10_c19 <= AA_c19(11);
   bh2012_wm29_11_c19 <= AA_c19(12);
   bh2012_wm28_9_c19 <= AA_c19(13);
   bh2012_wm27_9_c19 <= AA_c19(14);
   bh2012_wm26_9_c19 <= AA_c19(15);
   bh2012_wm25_10_c19 <= AA_c19(16);
   bh2012_wm24_9_c19 <= AA_c19(17);
   bh2012_wm23_9_c19 <= AA_c19(18);
   bh2012_wm22_9_c19 <= AA_c19(19);
   bh2012_wm21_10_c19 <= AA_c19(20);
   bh2012_wm20_8_c19 <= AA_c19(21);
   bh2012_wm19_9_c19 <= AA_c19(22);
   bh2012_wm18_9_c19 <= AA_c19(23);
   bh2012_wm17_8_c19 <= AA_c19(24);
   bh2012_wm16_8_c19 <= AA_c19(25);
   bh2012_wm15_7_c19 <= AA_c19(26);
   bh2012_wm14_5_c19 <= AA_c19(27);
   bh2012_wm13_5_c19 <= AA_c19(28);
   bh2012_wm12_5_c19 <= AA_c19(29);
   bh2012_wm11_3_c19 <= AA_c19(30);
   bh2012_wm10_2_c19 <= AA_c19(31);
   bh2012_wm9_2_c19 <= AA_c19(32);
   bh2012_wm8_1_c19 <= AA_c19(33);
   bh2012_wm7_0_c19 <= AA_c19(34);
   bh2012_wm6_0_c19 <= AA_c19(35);
   bh2012_wm5_0_c19 <= AA_c19(36);
   bh2012_wm4_0_c19 <= AA_c19(37);
   bh2012_wm3_0_c19 <= AA_c19(38);
   bh2012_wm2_0_c19 <= not AA_c19(39);

   -- Adding the constant bits 
   bh2012_wm42_5_c0 <= '1';
   bh2012_wm33_12_c0 <= '1';
   bh2012_wm32_11_c0 <= '1';
   bh2012_wm31_10_c0 <= '1';
   bh2012_wm30_11_c0 <= '1';
   bh2012_wm28_10_c0 <= '1';
   bh2012_wm27_10_c0 <= '1';
   bh2012_wm26_10_c0 <= '1';
   bh2012_wm24_10_c0 <= '1';
   bh2012_wm23_10_c0 <= '1';
   bh2012_wm22_10_c0 <= '1';
   bh2012_wm21_11_c0 <= '1';
   bh2012_wm19_10_c0 <= '1';
   bh2012_wm18_10_c0 <= '1';
   bh2012_wm14_6_c0 <= '1';
   bh2012_wm10_3_c0 <= '1';
   bh2012_wm7_1_c0 <= '1';
   bh2012_wm6_1_c0 <= '1';
   bh2012_wm5_1_c0 <= '1';
   bh2012_wm4_1_c0 <= '1';
   bh2012_wm3_1_c0 <= '1';
   bh2012_wm1_0_c0 <= '1';


   Compressor_23_3_Freq300_uid2256_bh2012_uid2257_In0_c22 <= "" & bh2012_wm52_0_c22 & bh2012_wm52_1_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2257_In1_c22 <= "" & bh2012_wm51_0_c22 & bh2012_wm51_1_c22;
   bh2012_wm52_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_c22(0);
   bh2012_wm51_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_c22(1);
   bh2012_wm50_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2257: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2257_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2257_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_copy2258_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2257_Out0_copy2258_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2259_In0_c22 <= "" & bh2012_wm50_0_c22 & bh2012_wm50_1_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2259_In1_c22 <= "" & bh2012_wm49_0_c22 & bh2012_wm49_1_c22;
   bh2012_wm50_3_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_c22(0);
   bh2012_wm49_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_c22(1);
   bh2012_wm48_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2259: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2259_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2259_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_copy2260_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2259_Out0_copy2260_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2261_In0_c22 <= "" & bh2012_wm48_0_c22 & bh2012_wm48_1_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2261_In1_c22 <= "" & bh2012_wm47_0_c22 & bh2012_wm47_1_c22;
   bh2012_wm48_3_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_c22(0);
   bh2012_wm47_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_c22(1);
   bh2012_wm46_2_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2261: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2261_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2261_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_copy2262_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2261_Out0_copy2262_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2265_In0_c22 <= "" & bh2012_wm46_0_c22 & bh2012_wm46_1_c22 & "0";
   bh2012_wm46_3_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_c22(0);
   bh2012_wm45_3_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2265: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2265_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_copy2266_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2265_Out0_copy2266_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2267_In0_c22 <= "" & bh2012_wm45_0_c22 & bh2012_wm45_1_c22 & bh2012_wm45_2_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2267_In1_c22 <= "" & bh2012_wm44_0_c22 & bh2012_wm44_1_c22;
   bh2012_wm45_4_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_c22(0);
   bh2012_wm44_3_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_c22(1);
   bh2012_wm43_4_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2267: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2267_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2267_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_copy2268_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2267_Out0_copy2268_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2269_In0_c22 <= "" & bh2012_wm43_0_c22 & bh2012_wm43_1_c22 & bh2012_wm43_2_c22;
   bh2012_wm43_5_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_c22(0);
   bh2012_wm42_6_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2269: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2269_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_copy2270_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2269_Out0_copy2270_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2273_In0_c22 <= "" & bh2012_wm42_0_c22 & bh2012_wm42_1_c22 & bh2012_wm42_2_c22 & bh2012_wm42_3_c22 & bh2012_wm42_4_c22 & bh2012_wm42_5_c22;
   bh2012_wm42_7_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_c22(0);
   bh2012_wm41_7_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_c22(1);
   bh2012_wm40_7_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2273: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2273_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_copy2274_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2273_Out0_copy2274_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2275_In0_c22 <= "" & bh2012_wm41_0_c22 & bh2012_wm41_1_c22 & bh2012_wm41_2_c22 & bh2012_wm41_3_c22 & bh2012_wm41_4_c22 & bh2012_wm41_5_c22;
   bh2012_wm41_8_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_c22(0);
   bh2012_wm40_8_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_c22(1);
   bh2012_wm39_9_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2275: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2275_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_copy2276_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2275_Out0_copy2276_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2277_In0_c22 <= "" & bh2012_wm40_0_c22 & bh2012_wm40_1_c22 & bh2012_wm40_2_c22 & bh2012_wm40_3_c22 & bh2012_wm40_4_c22 & bh2012_wm40_5_c22;
   bh2012_wm40_9_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_c22(0);
   bh2012_wm39_10_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_c22(1);
   bh2012_wm38_9_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2277: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2277_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_copy2278_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2277_Out0_copy2278_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2279_In0_c22 <= "" & bh2012_wm39_0_c22 & bh2012_wm39_1_c22 & bh2012_wm39_2_c22 & bh2012_wm39_3_c22 & bh2012_wm39_4_c22 & bh2012_wm39_5_c22;
   bh2012_wm39_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_c22(0);
   bh2012_wm38_10_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_c22(1);
   bh2012_wm37_10_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2279: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2279_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_copy2280_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2279_Out0_copy2280_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In0_c21 <= "" & bh2012_wm39_6_c21 & bh2012_wm39_7_c21 & bh2012_wm39_8_c21;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In1_c22 <= "" & bh2012_wm38_0_c22 & bh2012_wm38_1_c22;
   bh2012_wm39_12_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_c22(0);
   bh2012_wm38_11_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_c22(1);
   bh2012_wm37_11_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2281: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2281_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_copy2282_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2281_Out0_copy2282_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2283_In0_c21 <= "" & bh2012_wm38_2_c21 & bh2012_wm38_3_c21 & bh2012_wm38_4_c21 & bh2012_wm38_5_c21 & bh2012_wm38_6_c21 & bh2012_wm38_7_c21;
   bh2012_wm38_12_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_c21(0);
   bh2012_wm37_12_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_c21(1);
   bh2012_wm36_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2283: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2283_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_copy2284_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2283_Out0_copy2284_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2285_In0_c22 <= "" & bh2012_wm37_0_c22 & bh2012_wm37_1_c22 & bh2012_wm37_2_c22 & bh2012_wm37_3_c22 & bh2012_wm37_4_c22 & bh2012_wm37_5_c22;
   bh2012_wm37_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_c22(0);
   bh2012_wm36_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_c22(1);
   bh2012_wm35_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2285: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2285_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_copy2286_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2285_Out0_copy2286_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In0_c21 <= "" & bh2012_wm37_6_c21 & bh2012_wm37_7_c21 & bh2012_wm37_8_c21 & bh2012_wm37_9_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In1_c22 <= "" & bh2012_wm36_0_c22;
   bh2012_wm37_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_c22(0);
   bh2012_wm36_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_c22(1);
   bh2012_wm35_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2289: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2289_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_copy2290_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2289_Out0_copy2290_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2291_In0_c22 <= "" & bh2012_wm36_1_c22 & bh2012_wm36_2_c22 & bh2012_wm36_3_c22 & bh2012_wm36_4_c22 & bh2012_wm36_5_c22 & bh2012_wm36_6_c22;
   bh2012_wm36_14_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_c22(0);
   bh2012_wm35_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_c22(1);
   bh2012_wm34_10_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2291: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2291_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_copy2292_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2291_Out0_copy2292_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In0_c21 <= "" & bh2012_wm36_7_c21 & bh2012_wm36_8_c21 & bh2012_wm36_9_c21 & bh2012_wm36_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In1_c22 <= "" & bh2012_wm35_0_c22;
   bh2012_wm36_15_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_c22(0);
   bh2012_wm35_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_c22(1);
   bh2012_wm34_11_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2293: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2293_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_copy2294_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2293_Out0_copy2294_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2295_In0_c22 <= "" & bh2012_wm35_1_c22 & bh2012_wm35_2_c22 & bh2012_wm35_3_c22 & bh2012_wm35_4_c22 & bh2012_wm35_5_c22 & bh2012_wm35_6_c22;
   bh2012_wm35_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_c22(0);
   bh2012_wm34_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_c22(1);
   bh2012_wm33_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2295: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2295_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_copy2296_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2295_Out0_copy2296_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In0_c21 <= "" & bh2012_wm35_7_c21 & bh2012_wm35_8_c21 & bh2012_wm35_9_c21 & bh2012_wm35_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In1_c22 <= "" & bh2012_wm34_0_c22;
   bh2012_wm35_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_c22(0);
   bh2012_wm34_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_c22(1);
   bh2012_wm33_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2297: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2297_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_copy2298_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2297_Out0_copy2298_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2299_In0_c22 <= "" & bh2012_wm34_1_c22 & bh2012_wm34_2_c22 & bh2012_wm34_3_c22 & bh2012_wm34_4_c22 & bh2012_wm34_5_c22 & bh2012_wm34_6_c22;
   bh2012_wm34_14_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_c22(0);
   bh2012_wm33_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_c22(1);
   bh2012_wm32_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2299: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2299_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_copy2300_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2299_Out0_copy2300_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2301_In0_c21 <= "" & bh2012_wm34_7_c21 & bh2012_wm34_8_c21 & bh2012_wm34_9_c21;
   bh2012_wm34_15_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_c21(0);
   bh2012_wm33_16_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_c21(1);
   Compressor_3_2_Freq300_uid2264_uid2301: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2301_In0_c21,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_copy2302_c21);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2301_Out0_copy2302_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2303_In0_c22 <= "" & bh2012_wm33_8_c22 & bh2012_wm33_12_c22 & bh2012_wm33_11_c22 & bh2012_wm33_10_c22 & bh2012_wm33_9_c22 & bh2012_wm33_0_c22;
   bh2012_wm33_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_c22(0);
   bh2012_wm32_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_c22(1);
   bh2012_wm31_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2303: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2303_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_copy2304_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2303_Out0_copy2304_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2305_In0_c22 <= "" & bh2012_wm33_1_c22 & bh2012_wm33_2_c22 & bh2012_wm33_3_c22 & bh2012_wm33_4_c22 & bh2012_wm33_5_c22 & bh2012_wm33_6_c22;
   bh2012_wm33_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_c22(0);
   bh2012_wm32_14_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_c22(1);
   bh2012_wm31_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2305: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2305_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_copy2306_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2305_Out0_copy2306_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2307_In0_c22 <= "" & bh2012_wm32_0_c22 & bh2012_wm32_1_c22 & bh2012_wm32_2_c22 & bh2012_wm32_3_c22 & bh2012_wm32_4_c22 & bh2012_wm32_5_c22;
   bh2012_wm32_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_c22(0);
   bh2012_wm31_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_c22(1);
   bh2012_wm30_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2307: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2307_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_copy2308_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2307_Out0_copy2308_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2309_In0_c21 <= "" & bh2012_wm32_6_c21 & bh2012_wm32_7_c21 & bh2012_wm32_8_c21 & bh2012_wm32_9_c21 & bh2012_wm32_10_c21 & bh2012_wm32_11_c21;
   bh2012_wm32_16_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_c21(0);
   bh2012_wm31_14_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_c21(1);
   bh2012_wm30_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2309: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2309_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_copy2310_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2309_Out0_copy2310_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2311_In0_c22 <= "" & bh2012_wm31_0_c22 & bh2012_wm31_1_c22 & bh2012_wm31_2_c22 & bh2012_wm31_3_c22 & bh2012_wm31_4_c22 & bh2012_wm31_5_c22;
   bh2012_wm31_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_c22(0);
   bh2012_wm30_14_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_c22(1);
   bh2012_wm29_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2311: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2311_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_copy2312_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2311_Out0_copy2312_c22; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid2314_bh2012_uid2315_In0_c21 <= "" & bh2012_wm31_6_c21 & bh2012_wm31_7_c21 & bh2012_wm31_8_c21 & bh2012_wm31_9_c21 & bh2012_wm31_10_c21;
   bh2012_wm31_16_c21 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_c21(0);
   bh2012_wm30_15_c21 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_c21(1);
   bh2012_wm29_13_c21 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_c21(2);
   Compressor_5_3_Freq300_uid2314_uid2315: Compressor_5_3_Freq300_uid2314
      port map ( X0 => Compressor_5_3_Freq300_uid2314_bh2012_uid2315_In0_c21,
                 R => Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_copy2316_c21);
   Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_c21 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2315_Out0_copy2316_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2317_In0_c22 <= "" & bh2012_wm30_0_c22 & bh2012_wm30_1_c22 & bh2012_wm30_2_c22 & bh2012_wm30_3_c22 & bh2012_wm30_4_c22 & bh2012_wm30_5_c22;
   bh2012_wm30_16_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_c22(0);
   bh2012_wm29_14_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_c22(1);
   bh2012_wm28_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2317: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2317_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_copy2318_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2317_Out0_copy2318_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2319_In0_c21 <= "" & bh2012_wm30_8_c21 & bh2012_wm30_11_c21 & bh2012_wm30_10_c21 & bh2012_wm30_9_c21 & bh2012_wm30_7_c21 & bh2012_wm30_6_c21;
   bh2012_wm30_17_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_c21(0);
   bh2012_wm29_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_c21(1);
   bh2012_wm28_12_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2319: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2319_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_copy2320_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2319_Out0_copy2320_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2321_In0_c22 <= "" & bh2012_wm29_0_c22 & bh2012_wm29_1_c22 & bh2012_wm29_2_c22 & bh2012_wm29_3_c22 & bh2012_wm29_4_c22 & bh2012_wm29_5_c22;
   bh2012_wm29_16_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_c22(0);
   bh2012_wm28_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_c22(1);
   bh2012_wm27_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2321: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2321_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_copy2322_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2321_Out0_copy2322_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2323_In0_c21 <= "" & bh2012_wm29_8_c21 & bh2012_wm29_11_c21 & bh2012_wm29_10_c21 & bh2012_wm29_9_c21 & bh2012_wm29_7_c21 & bh2012_wm29_6_c21;
   bh2012_wm29_17_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_c21(0);
   bh2012_wm28_14_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_c21(1);
   bh2012_wm27_12_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2323: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2323_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_copy2324_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2323_Out0_copy2324_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2325_In0_c22 <= "" & bh2012_wm28_0_c22 & bh2012_wm28_1_c22 & bh2012_wm28_2_c22 & bh2012_wm28_3_c22 & bh2012_wm28_4_c22 & bh2012_wm28_5_c22;
   bh2012_wm28_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_c22(0);
   bh2012_wm27_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_c22(1);
   bh2012_wm26_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2325: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2325_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_copy2326_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2325_Out0_copy2326_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In0_c21 <= "" & bh2012_wm28_6_c21 & bh2012_wm28_7_c21 & bh2012_wm28_8_c21 & bh2012_wm28_9_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In1_c22 <= "" & bh2012_wm27_0_c22;
   bh2012_wm28_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_c22(0);
   bh2012_wm27_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_c22(1);
   bh2012_wm26_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2327: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2327_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_copy2328_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2327_Out0_copy2328_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2329_In0_c21 <= "" & bh2012_wm27_1_c21 & bh2012_wm27_2_c21 & bh2012_wm27_3_c21 & bh2012_wm27_4_c21 & bh2012_wm27_5_c21 & bh2012_wm27_6_c21;
   bh2012_wm27_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_c21(0);
   bh2012_wm26_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_c21(1);
   bh2012_wm25_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2329: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2329_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_copy2330_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2329_Out0_copy2330_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In0_c21 <= "" & bh2012_wm27_7_c21 & bh2012_wm27_8_c21 & bh2012_wm27_9_c21 & bh2012_wm27_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In1_c22 <= "" & bh2012_wm26_0_c22;
   bh2012_wm27_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_c22(0);
   bh2012_wm26_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_c22(1);
   bh2012_wm25_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2331: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2331_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_copy2332_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2331_Out0_copy2332_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2333_In0_c21 <= "" & bh2012_wm26_1_c21 & bh2012_wm26_2_c21 & bh2012_wm26_3_c21 & bh2012_wm26_4_c21 & bh2012_wm26_5_c21 & bh2012_wm26_6_c21;
   bh2012_wm26_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_c21(0);
   bh2012_wm25_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_c21(1);
   bh2012_wm24_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2333: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2333_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_copy2334_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2333_Out0_copy2334_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In0_c21 <= "" & bh2012_wm26_7_c21 & bh2012_wm26_8_c21 & bh2012_wm26_9_c21 & bh2012_wm26_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In1_c22 <= "" & bh2012_wm25_0_c22;
   bh2012_wm26_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_c22(0);
   bh2012_wm25_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_c22(1);
   bh2012_wm24_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2335: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2335_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_copy2336_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2335_Out0_copy2336_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2337_In0_c21 <= "" & bh2012_wm25_1_c21 & bh2012_wm25_2_c21 & bh2012_wm25_3_c21 & bh2012_wm25_4_c21 & bh2012_wm25_5_c21 & bh2012_wm25_6_c21;
   bh2012_wm25_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_c21(0);
   bh2012_wm24_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_c21(1);
   bh2012_wm23_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2337: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2337_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_copy2338_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2337_Out0_copy2338_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In0_c21 <= "" & bh2012_wm25_7_c21 & bh2012_wm25_8_c21 & bh2012_wm25_9_c21 & bh2012_wm25_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In1_c22 <= "" & bh2012_wm24_0_c22;
   bh2012_wm25_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_c22(0);
   bh2012_wm24_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_c22(1);
   bh2012_wm23_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2339: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2339_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_copy2340_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2339_Out0_copy2340_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2341_In0_c21 <= "" & bh2012_wm24_1_c21 & bh2012_wm24_2_c21 & bh2012_wm24_3_c21 & bh2012_wm24_4_c21 & bh2012_wm24_5_c21 & bh2012_wm24_6_c21;
   bh2012_wm24_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_c21(0);
   bh2012_wm23_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_c21(1);
   bh2012_wm22_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2341: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2341_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_copy2342_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2341_Out0_copy2342_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In0_c21 <= "" & bh2012_wm24_7_c21 & bh2012_wm24_8_c21 & bh2012_wm24_9_c21 & bh2012_wm24_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In1_c22 <= "" & bh2012_wm23_0_c22;
   bh2012_wm24_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_c22(0);
   bh2012_wm23_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_c22(1);
   bh2012_wm22_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2343: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2343_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_copy2344_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2343_Out0_copy2344_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2345_In0_c21 <= "" & bh2012_wm23_1_c21 & bh2012_wm23_2_c21 & bh2012_wm23_3_c21 & bh2012_wm23_4_c21 & bh2012_wm23_5_c21 & bh2012_wm23_6_c21;
   bh2012_wm23_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_c21(0);
   bh2012_wm22_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_c21(1);
   bh2012_wm21_12_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2345: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2345_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_copy2346_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2345_Out0_copy2346_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In0_c21 <= "" & bh2012_wm23_7_c21 & bh2012_wm23_8_c21 & bh2012_wm23_9_c21 & bh2012_wm23_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In1_c22 <= "" & bh2012_wm22_0_c22;
   bh2012_wm23_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_c22(0);
   bh2012_wm22_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_c22(1);
   bh2012_wm21_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2347: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2347_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_copy2348_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2347_Out0_copy2348_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2349_In0_c21 <= "" & bh2012_wm22_1_c21 & bh2012_wm22_2_c21 & bh2012_wm22_3_c21 & bh2012_wm22_4_c21 & bh2012_wm22_5_c21 & bh2012_wm22_6_c21;
   bh2012_wm22_15_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_c21(0);
   bh2012_wm21_14_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_c21(1);
   bh2012_wm20_9_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2349: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2349_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_copy2350_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2349_Out0_copy2350_c21; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2351_In0_c21 <= "" & bh2012_wm22_7_c21 & bh2012_wm22_8_c21 & bh2012_wm22_9_c21;
   bh2012_wm22_16_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_c21(0);
   bh2012_wm21_15_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_c21(1);
   Compressor_3_2_Freq300_uid2264_uid2351: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2351_In0_c21,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_copy2352_c21);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2351_Out0_copy2352_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2353_In0_c22 <= "" & bh2012_wm21_0_c22 & bh2012_wm21_1_c22 & bh2012_wm21_2_c22 & bh2012_wm21_3_c22 & bh2012_wm21_4_c22 & bh2012_wm21_5_c22;
   bh2012_wm21_16_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_c22(0);
   bh2012_wm20_10_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_c22(1);
   bh2012_wm19_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2353: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2353_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_copy2354_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2353_Out0_copy2354_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2355_In0_c21 <= "" & bh2012_wm21_8_c21 & bh2012_wm21_11_c21 & bh2012_wm21_10_c21 & bh2012_wm21_9_c21 & bh2012_wm21_7_c21 & bh2012_wm21_6_c21;
   bh2012_wm21_17_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_c21(0);
   bh2012_wm20_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_c21(1);
   bh2012_wm19_12_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2355: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2355_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_copy2356_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2355_Out0_copy2356_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2357_In0_c22 <= "" & bh2012_wm20_0_c22 & bh2012_wm20_1_c22 & bh2012_wm20_2_c22 & bh2012_wm20_3_c22 & bh2012_wm20_4_c22 & bh2012_wm20_5_c22;
   bh2012_wm20_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_c22(0);
   bh2012_wm19_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_c22(1);
   bh2012_wm18_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2357: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2357_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_copy2358_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2357_Out0_copy2358_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2359_In0_c21 <= "" & bh2012_wm20_6_c21 & bh2012_wm20_7_c21 & bh2012_wm20_8_c21;
   bh2012_wm20_13_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_c21(0);
   bh2012_wm19_14_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_c21(1);
   Compressor_3_2_Freq300_uid2264_uid2359: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2359_In0_c21,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_copy2360_c21);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2359_Out0_copy2360_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2361_In0_c22 <= "" & bh2012_wm19_0_c22 & bh2012_wm19_1_c22 & bh2012_wm19_2_c22 & bh2012_wm19_3_c22 & bh2012_wm19_4_c22 & bh2012_wm19_5_c22;
   bh2012_wm19_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_c22(0);
   bh2012_wm18_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_c22(1);
   bh2012_wm17_9_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2361: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2361_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_copy2362_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2361_Out0_copy2362_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In0_c21 <= "" & bh2012_wm19_6_c21 & bh2012_wm19_7_c21 & bh2012_wm19_8_c21 & bh2012_wm19_9_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In1_c22 <= "" & bh2012_wm18_0_c22;
   bh2012_wm19_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_c22(0);
   bh2012_wm18_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_c22(1);
   bh2012_wm17_10_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2363: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2363_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_copy2364_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2363_Out0_copy2364_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2365_In0_c21 <= "" & bh2012_wm18_1_c21 & bh2012_wm18_2_c21 & bh2012_wm18_3_c21 & bh2012_wm18_4_c21 & bh2012_wm18_5_c21 & bh2012_wm18_6_c21;
   bh2012_wm18_14_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_c21(0);
   bh2012_wm17_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_c21(1);
   bh2012_wm16_9_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2365: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2365_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_copy2366_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2365_Out0_copy2366_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In0_c21 <= "" & bh2012_wm18_7_c21 & bh2012_wm18_8_c21 & bh2012_wm18_9_c21 & bh2012_wm18_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c0 <= "" & "0";
   bh2012_wm18_15_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_c21(0);
   bh2012_wm17_12_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_c21(1);
   bh2012_wm16_10_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_c21(2);
   Compressor_14_3_Freq300_uid2288_uid2367: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In0_c21,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2367_In1_c21,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_copy2368_c21);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2367_Out0_copy2368_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2369_In0_c22 <= "" & bh2012_wm17_0_c22 & bh2012_wm17_1_c22 & bh2012_wm17_2_c22 & bh2012_wm17_3_c22 & bh2012_wm17_4_c22 & bh2012_wm17_5_c22;
   bh2012_wm17_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_c22(0);
   bh2012_wm16_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_c22(1);
   bh2012_wm15_8_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2369: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2369_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_copy2370_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2369_Out0_copy2370_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2371_In0_c21 <= "" & bh2012_wm17_6_c21 & bh2012_wm17_7_c21 & bh2012_wm17_8_c21;
   bh2012_wm17_14_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_c21(0);
   bh2012_wm16_12_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_c21(1);
   Compressor_3_2_Freq300_uid2264_uid2371: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2371_In0_c21,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_copy2372_c21);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_c21 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2371_Out0_copy2372_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2373_In0_c21 <= "" & bh2012_wm16_0_c21 & bh2012_wm16_1_c21 & bh2012_wm16_2_c21 & bh2012_wm16_3_c21 & bh2012_wm16_4_c21 & bh2012_wm16_5_c21;
   bh2012_wm16_13_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_c21(0);
   bh2012_wm15_9_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_c21(1);
   bh2012_wm14_7_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2373: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2373_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_copy2374_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2373_Out0_copy2374_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2375_In0_c21 <= "" & bh2012_wm16_6_c21 & bh2012_wm16_7_c21 & bh2012_wm16_8_c21;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2375_In1_c21 <= "" & bh2012_wm15_0_c21 & bh2012_wm15_1_c21;
   bh2012_wm16_14_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_c21(0);
   bh2012_wm15_10_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_c21(1);
   bh2012_wm14_8_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_c21(2);
   Compressor_23_3_Freq300_uid2256_uid2375: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2375_In0_c21,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2375_In1_c21,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_copy2376_c21);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2375_Out0_copy2376_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2377_In0_c21 <= "" & bh2012_wm15_2_c21 & bh2012_wm15_3_c21 & bh2012_wm15_4_c21 & bh2012_wm15_5_c21 & bh2012_wm15_6_c21 & bh2012_wm15_7_c21;
   bh2012_wm15_11_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_c21(0);
   bh2012_wm14_9_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_c21(1);
   bh2012_wm13_6_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2377: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2377_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_copy2378_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2377_Out0_copy2378_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2379_In0_c21 <= "" & bh2012_wm14_0_c21 & bh2012_wm14_1_c21 & bh2012_wm14_2_c21 & bh2012_wm14_3_c21 & bh2012_wm14_4_c21 & bh2012_wm14_5_c21;
   bh2012_wm14_10_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_c21(0);
   bh2012_wm13_7_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_c21(1);
   bh2012_wm12_6_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2379: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2379_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_copy2380_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2379_Out0_copy2380_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2381_In0_c21 <= "" & bh2012_wm13_0_c21 & bh2012_wm13_1_c21 & bh2012_wm13_2_c21 & bh2012_wm13_3_c21 & bh2012_wm13_4_c21 & bh2012_wm13_5_c21;
   bh2012_wm13_8_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_c21(0);
   bh2012_wm12_7_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_c21(1);
   bh2012_wm11_4_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2381: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2381_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_copy2382_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2381_Out0_copy2382_c21; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2383_In0_c21 <= "" & bh2012_wm12_0_c21 & bh2012_wm12_1_c21 & bh2012_wm12_2_c21 & bh2012_wm12_3_c21 & bh2012_wm12_4_c21 & bh2012_wm12_5_c21;
   bh2012_wm12_8_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_c21(0);
   bh2012_wm11_5_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_c21(1);
   bh2012_wm10_4_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_c21(2);
   Compressor_6_3_Freq300_uid2272_uid2383: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2383_In0_c21,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_copy2384_c21);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_c21 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2383_Out0_copy2384_c21; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2385_In0_c21 <= "" & bh2012_wm11_0_c21 & bh2012_wm11_1_c21 & bh2012_wm11_2_c21 & bh2012_wm11_3_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2385_In1_c21 <= "" & bh2012_wm10_0_c21;
   bh2012_wm11_6_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_c21(0);
   bh2012_wm10_5_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_c21(1);
   bh2012_wm9_3_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_c21(2);
   Compressor_14_3_Freq300_uid2288_uid2385: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2385_In0_c21,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2385_In1_c21,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_copy2386_c21);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_c21 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2385_Out0_copy2386_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2387_In0_c21 <= "" & bh2012_wm10_1_c21 & bh2012_wm10_2_c21 & bh2012_wm10_3_c21;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2387_In1_c21 <= "" & bh2012_wm9_0_c21 & bh2012_wm9_1_c21;
   bh2012_wm10_6_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_c21(0);
   bh2012_wm9_4_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_c21(1);
   bh2012_wm8_2_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_c21(2);
   Compressor_23_3_Freq300_uid2256_uid2387: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2387_In0_c21,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2387_In1_c21,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_copy2388_c21);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2387_Out0_copy2388_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In0_c21 <= "" & bh2012_wm8_0_c21 & bh2012_wm8_1_c21 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c19 <= "" & bh2012_wm7_0_c19 & bh2012_wm7_1_c19;
   bh2012_wm8_3_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_c21(0);
   bh2012_wm7_2_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_c21(1);
   bh2012_wm6_2_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_c21(2);
   Compressor_23_3_Freq300_uid2256_uid2389: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In0_c21,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2389_In1_c21,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_copy2390_c21);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_c21 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2389_Out0_copy2390_c21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2391_In0_c19 <= "" & bh2012_wm6_0_c19 & bh2012_wm6_1_c19 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2391_In1_c19 <= "" & bh2012_wm5_0_c19 & bh2012_wm5_1_c19;
   bh2012_wm6_3_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_c19(0);
   bh2012_wm5_2_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_c19(1);
   bh2012_wm4_2_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_c19(2);
   Compressor_23_3_Freq300_uid2256_uid2391: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2391_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2391_In1_c19,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_copy2392_c19);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2391_Out0_copy2392_c19; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2393_In0_c19 <= "" & bh2012_wm4_0_c19 & bh2012_wm4_1_c19 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2393_In1_c19 <= "" & bh2012_wm3_0_c19 & bh2012_wm3_1_c19;
   bh2012_wm4_3_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_c19(0);
   bh2012_wm3_2_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_c19(1);
   bh2012_wm2_1_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_c19(2);
   Compressor_23_3_Freq300_uid2256_uid2393: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2393_In0_c19,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2393_In1_c19,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_copy2394_c19);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_c19 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2393_Out0_copy2394_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2395_In0_c22 <= "" & bh2012_wm50_2_c22 & bh2012_wm50_3_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2395_In1_c22 <= "" & bh2012_wm49_2_c22;
   bh2012_wm50_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_c22(0);
   bh2012_wm49_3_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_c22(1);
   bh2012_wm48_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2395: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2395_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2395_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_copy2396_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2395_Out0_copy2396_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2397_In0_c22 <= "" & bh2012_wm48_2_c22 & bh2012_wm48_3_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2397_In1_c22 <= "" & bh2012_wm47_2_c22;
   bh2012_wm48_5_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_c22(0);
   bh2012_wm47_3_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_c22(1);
   bh2012_wm46_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2397: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2397_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2397_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_copy2398_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2397_Out0_copy2398_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2399_In0_c22 <= "" & bh2012_wm46_2_c22 & bh2012_wm46_3_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2399_In1_c22 <= "" & bh2012_wm45_3_c22 & bh2012_wm45_4_c22;
   bh2012_wm46_5_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_c22(0);
   bh2012_wm45_5_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_c22(1);
   bh2012_wm44_4_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2399: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2399_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2399_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_copy2400_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2399_Out0_copy2400_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2401_In0_c22 <= "" & bh2012_wm44_2_c22 & bh2012_wm44_3_c22 & "0";
   bh2012_wm44_5_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_c22(0);
   bh2012_wm43_6_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2401: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2401_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_copy2402_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2401_Out0_copy2402_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2403_In0_c22 <= "" & bh2012_wm43_3_c22 & bh2012_wm43_4_c22 & bh2012_wm43_5_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2403_In1_c22 <= "" & bh2012_wm42_6_c22 & bh2012_wm42_7_c22;
   bh2012_wm43_7_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_c22(0);
   bh2012_wm42_8_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_c22(1);
   bh2012_wm41_9_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2403: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2403_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2403_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_copy2404_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2403_Out0_copy2404_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2405_In0_c22 <= "" & bh2012_wm41_6_c22 & bh2012_wm41_7_c22 & bh2012_wm41_8_c22;
   bh2012_wm41_10_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_c22(0);
   bh2012_wm40_10_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2405: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2405_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_copy2406_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2405_Out0_copy2406_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2407_In0_c22 <= "" & bh2012_wm40_6_c22 & bh2012_wm40_7_c22 & bh2012_wm40_8_c22 & bh2012_wm40_9_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2407_In1_c22 <= "" & bh2012_wm39_9_c22;
   bh2012_wm40_11_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_c22(0);
   bh2012_wm39_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_c22(1);
   bh2012_wm38_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2407: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2407_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2407_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_copy2408_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2407_Out0_copy2408_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2409_In0_c22 <= "" & bh2012_wm39_10_c22 & bh2012_wm39_11_c22 & bh2012_wm39_12_c22;
   bh2012_wm39_14_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_c22(0);
   bh2012_wm38_14_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2409: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2409_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_copy2410_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2409_Out0_copy2410_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2411_In0_c22 <= "" & bh2012_wm38_8_c22 & bh2012_wm38_9_c22 & bh2012_wm38_10_c22 & bh2012_wm38_11_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2411_In1_c22 <= "" & bh2012_wm37_10_c22;
   bh2012_wm38_15_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_c22(0);
   bh2012_wm37_15_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_c22(1);
   bh2012_wm36_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2411: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2411_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2411_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_copy2412_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2411_Out0_copy2412_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In0_c22 <= "" & bh2012_wm37_11_c22 & bh2012_wm37_12_c22 & bh2012_wm37_13_c22 & bh2012_wm37_14_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In1_c21 <= "" & bh2012_wm36_11_c21;
   bh2012_wm37_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_c22(0);
   bh2012_wm36_17_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_c22(1);
   bh2012_wm35_17_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2413: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2413_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_copy2414_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2413_Out0_copy2414_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2415_In0_c22 <= "" & bh2012_wm36_12_c22 & bh2012_wm36_13_c22 & bh2012_wm36_14_c22;
   bh2012_wm36_18_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_c22(0);
   bh2012_wm35_18_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2415: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2415_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_copy2416_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2415_Out0_copy2416_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2417_In0_c22 <= "" & bh2012_wm35_11_c22 & bh2012_wm35_12_c22 & bh2012_wm35_13_c22 & bh2012_wm35_14_c22 & bh2012_wm35_15_c22 & bh2012_wm35_16_c22;
   bh2012_wm35_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_c22(0);
   bh2012_wm34_16_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_c22(1);
   bh2012_wm33_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2417: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2417_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_copy2418_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2417_Out0_copy2418_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2419_In0_c22 <= "" & bh2012_wm34_10_c22 & bh2012_wm34_11_c22 & bh2012_wm34_12_c22 & bh2012_wm34_13_c22 & bh2012_wm34_14_c22 & bh2012_wm34_15_c22;
   bh2012_wm34_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_c22(0);
   bh2012_wm33_20_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_c22(1);
   bh2012_wm32_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2419: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2419_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_copy2420_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2419_Out0_copy2420_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2421_In0_c22 <= "" & bh2012_wm33_17_c22 & bh2012_wm33_7_c22 & bh2012_wm33_13_c22 & bh2012_wm33_14_c22 & bh2012_wm33_15_c22 & bh2012_wm33_16_c22;
   bh2012_wm33_21_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_c22(0);
   bh2012_wm32_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_c22(1);
   bh2012_wm31_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2421: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2421_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_copy2422_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2421_Out0_copy2422_c22; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid2314_bh2012_uid2423_In0_c22 <= "" & bh2012_wm32_12_c22 & bh2012_wm32_13_c22 & bh2012_wm32_14_c22 & bh2012_wm32_15_c22 & bh2012_wm32_16_c22;
   bh2012_wm32_19_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_c22(0);
   bh2012_wm31_18_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_c22(1);
   bh2012_wm30_18_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_c22(2);
   Compressor_5_3_Freq300_uid2314_uid2423: Compressor_5_3_Freq300_uid2314
      port map ( X0 => Compressor_5_3_Freq300_uid2314_bh2012_uid2423_In0_c22,
                 R => Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_copy2424_c22);
   Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2423_Out0_copy2424_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2425_In0_c22 <= "" & bh2012_wm31_11_c22 & bh2012_wm31_12_c22 & bh2012_wm31_13_c22 & bh2012_wm31_14_c22 & bh2012_wm31_15_c22 & bh2012_wm31_16_c22;
   bh2012_wm31_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_c22(0);
   bh2012_wm30_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_c22(1);
   bh2012_wm29_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2425: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2425_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_copy2426_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2425_Out0_copy2426_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2427_In0_c22 <= "" & bh2012_wm30_16_c22 & bh2012_wm30_15_c22 & bh2012_wm30_14_c22 & bh2012_wm30_13_c22 & bh2012_wm30_12_c22 & bh2012_wm30_17_c22;
   bh2012_wm30_20_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_c22(0);
   bh2012_wm29_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_c22(1);
   bh2012_wm28_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2427: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2427_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_copy2428_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2427_Out0_copy2428_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2429_In0_c22 <= "" & bh2012_wm29_16_c22 & bh2012_wm29_15_c22 & bh2012_wm29_14_c22 & bh2012_wm29_13_c22 & bh2012_wm29_12_c22 & bh2012_wm29_17_c22;
   bh2012_wm29_20_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_c22(0);
   bh2012_wm28_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_c22(1);
   bh2012_wm27_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2429: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2429_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_copy2430_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2429_Out0_copy2430_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2431_In0_c22 <= "" & bh2012_wm28_10_c22 & bh2012_wm28_11_c22 & bh2012_wm28_12_c22 & bh2012_wm28_13_c22 & bh2012_wm28_14_c22 & bh2012_wm28_15_c22;
   bh2012_wm28_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_c22(0);
   bh2012_wm27_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_c22(1);
   bh2012_wm26_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2431: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2431_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_copy2432_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2431_Out0_copy2432_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2433_In0_c22 <= "" & bh2012_wm27_11_c22 & bh2012_wm27_12_c22 & bh2012_wm27_13_c22 & bh2012_wm27_14_c22 & bh2012_wm27_15_c22 & bh2012_wm27_16_c22;
   bh2012_wm27_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_c22(0);
   bh2012_wm26_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_c22(1);
   bh2012_wm25_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2433: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2433_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_copy2434_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2433_Out0_copy2434_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2435_In0_c22 <= "" & bh2012_wm26_11_c22 & bh2012_wm26_12_c22 & bh2012_wm26_13_c22 & bh2012_wm26_14_c22 & bh2012_wm26_15_c22 & bh2012_wm26_16_c22;
   bh2012_wm26_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_c22(0);
   bh2012_wm25_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_c22(1);
   bh2012_wm24_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2435: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2435_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_copy2436_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2435_Out0_copy2436_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2437_In0_c22 <= "" & bh2012_wm25_11_c22 & bh2012_wm25_12_c22 & bh2012_wm25_13_c22 & bh2012_wm25_14_c22 & bh2012_wm25_15_c22 & bh2012_wm25_16_c22;
   bh2012_wm25_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_c22(0);
   bh2012_wm24_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_c22(1);
   bh2012_wm23_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2437: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2437_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_copy2438_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2437_Out0_copy2438_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2439_In0_c22 <= "" & bh2012_wm24_11_c22 & bh2012_wm24_12_c22 & bh2012_wm24_13_c22 & bh2012_wm24_14_c22 & bh2012_wm24_15_c22 & bh2012_wm24_16_c22;
   bh2012_wm24_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_c22(0);
   bh2012_wm23_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_c22(1);
   bh2012_wm22_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2439: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2439_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_copy2440_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2439_Out0_copy2440_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2441_In0_c22 <= "" & bh2012_wm23_11_c22 & bh2012_wm23_12_c22 & bh2012_wm23_13_c22 & bh2012_wm23_14_c22 & bh2012_wm23_15_c22 & bh2012_wm23_16_c22;
   bh2012_wm23_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_c22(0);
   bh2012_wm22_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_c22(1);
   bh2012_wm21_18_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2441: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2441_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_copy2442_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2441_Out0_copy2442_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2443_In0_c22 <= "" & bh2012_wm22_10_c22 & bh2012_wm22_11_c22 & bh2012_wm22_12_c22 & bh2012_wm22_13_c22 & bh2012_wm22_14_c22 & bh2012_wm22_15_c22;
   bh2012_wm22_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_c22(0);
   bh2012_wm21_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_c22(1);
   bh2012_wm20_14_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2443: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2443_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_copy2444_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2443_Out0_copy2444_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2445_In0_c22 <= "" & bh2012_wm21_16_c22 & bh2012_wm21_15_c22 & bh2012_wm21_14_c22 & bh2012_wm21_13_c22 & bh2012_wm21_12_c22 & bh2012_wm21_17_c22;
   bh2012_wm21_20_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_c22(0);
   bh2012_wm20_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_c22(1);
   bh2012_wm19_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2445: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2445_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_copy2446_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2445_Out0_copy2446_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In0_c22 <= "" & bh2012_wm20_9_c22 & bh2012_wm20_10_c22 & bh2012_wm20_11_c22 & bh2012_wm20_12_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c0 <= "" & bh2012_wm19_10_c0;
   bh2012_wm20_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_c22(0);
   bh2012_wm19_18_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_c22(1);
   bh2012_wm18_16_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2447: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2447_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_copy2448_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2447_Out0_copy2448_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2449_In0_c22 <= "" & bh2012_wm19_11_c22 & bh2012_wm19_12_c22 & bh2012_wm19_13_c22 & bh2012_wm19_14_c22 & bh2012_wm19_15_c22 & bh2012_wm19_16_c22;
   bh2012_wm19_19_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_c22(0);
   bh2012_wm18_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_c22(1);
   bh2012_wm17_15_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2449: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2449_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_copy2450_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2449_Out0_copy2450_c22; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid2314_bh2012_uid2451_In0_c22 <= "" & bh2012_wm18_11_c22 & bh2012_wm18_12_c22 & bh2012_wm18_13_c22 & bh2012_wm18_14_c22 & bh2012_wm18_15_c22;
   bh2012_wm18_18_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_c22(0);
   bh2012_wm17_16_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_c22(1);
   bh2012_wm16_15_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_c22(2);
   Compressor_5_3_Freq300_uid2314_uid2451: Compressor_5_3_Freq300_uid2314
      port map ( X0 => Compressor_5_3_Freq300_uid2314_bh2012_uid2451_In0_c22,
                 R => Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_copy2452_c22);
   Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_c22 <= Compressor_5_3_Freq300_uid2314_bh2012_uid2451_Out0_copy2452_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2453_In0_c22 <= "" & bh2012_wm17_9_c22 & bh2012_wm17_10_c22 & bh2012_wm17_11_c22 & bh2012_wm17_12_c22 & bh2012_wm17_13_c22 & bh2012_wm17_14_c22;
   bh2012_wm17_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_c22(0);
   bh2012_wm16_16_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_c22(1);
   bh2012_wm15_12_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2453: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2453_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_copy2454_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2453_Out0_copy2454_c22; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2272_bh2012_uid2455_In0_c22 <= "" & bh2012_wm16_9_c22 & bh2012_wm16_10_c22 & bh2012_wm16_11_c22 & bh2012_wm16_12_c22 & bh2012_wm16_13_c22 & bh2012_wm16_14_c22;
   bh2012_wm16_17_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_c22(0);
   bh2012_wm15_13_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_c22(1);
   bh2012_wm14_11_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_c22(2);
   Compressor_6_3_Freq300_uid2272_uid2455: Compressor_6_3_Freq300_uid2272
      port map ( X0 => Compressor_6_3_Freq300_uid2272_bh2012_uid2455_In0_c22,
                 R => Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_copy2456_c22);
   Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_c22 <= Compressor_6_3_Freq300_uid2272_bh2012_uid2455_Out0_copy2456_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In0_c22 <= "" & bh2012_wm15_8_c22 & bh2012_wm15_9_c22 & bh2012_wm15_10_c22 & bh2012_wm15_11_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c0 <= "" & bh2012_wm14_6_c0;
   bh2012_wm15_14_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_c22(0);
   bh2012_wm14_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_c22(1);
   bh2012_wm13_9_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2457: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2457_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_copy2458_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2457_Out0_copy2458_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In0_c21 <= "" & bh2012_wm14_7_c21 & bh2012_wm14_8_c21 & bh2012_wm14_9_c21 & bh2012_wm14_10_c21;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c0 <= "" & "0";
   bh2012_wm14_13_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_c22(0);
   bh2012_wm13_10_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_c22(1);
   bh2012_wm12_9_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2459: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In0_c21,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2459_In1_c21,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_copy2460_c21);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2459_Out0_copy2460_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2461_In0_c21 <= "" & bh2012_wm13_6_c21 & bh2012_wm13_7_c21 & bh2012_wm13_8_c21;
   bh2012_wm13_11_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_c22(0);
   bh2012_wm12_10_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2461: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2461_In0_c21,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_copy2462_c21);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2461_Out0_copy2462_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2463_In0_c21 <= "" & bh2012_wm12_6_c21 & bh2012_wm12_7_c21 & bh2012_wm12_8_c21;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2463_In1_c21 <= "" & bh2012_wm11_4_c21 & bh2012_wm11_5_c21;
   bh2012_wm12_11_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_c22(0);
   bh2012_wm11_7_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_c22(1);
   bh2012_wm10_7_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2463: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2463_In0_c21,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2463_In1_c21,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_copy2464_c21);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2463_Out0_copy2464_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2465_In0_c21 <= "" & bh2012_wm10_4_c21 & bh2012_wm10_5_c21 & bh2012_wm10_6_c21;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2465_In1_c21 <= "" & bh2012_wm9_2_c21 & bh2012_wm9_3_c21;
   bh2012_wm10_8_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_c22(0);
   bh2012_wm9_5_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_c22(1);
   bh2012_wm8_4_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2465: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2465_In0_c21,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2465_In1_c21,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_copy2466_c21);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2465_Out0_copy2466_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2467_In0_c21 <= "" & bh2012_wm8_2_c21 & bh2012_wm8_3_c21 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2467_In1_c21 <= "" & bh2012_wm7_2_c21;
   bh2012_wm8_5_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_c22(0);
   bh2012_wm7_3_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_c22(1);
   bh2012_wm6_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2467: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2467_In0_c21,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2467_In1_c21,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_copy2468_c21);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2467_Out0_copy2468_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In0_c21 <= "" & bh2012_wm6_2_c21 & bh2012_wm6_3_c21 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c19 <= "" & bh2012_wm5_2_c19;
   bh2012_wm6_5_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_c22(0);
   bh2012_wm5_3_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_c22(1);
   bh2012_wm4_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2469: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In0_c21,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2469_In1_c21,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_copy2470_c21);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2469_Out0_copy2470_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2471_In0_c19 <= "" & bh2012_wm4_2_c19 & bh2012_wm4_3_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2471_In1_c19 <= "" & bh2012_wm3_2_c19;
   bh2012_wm4_5_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_c19(0);
   bh2012_wm3_3_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_c19(1);
   bh2012_wm2_2_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_c19(2);
   Compressor_14_3_Freq300_uid2288_uid2471: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2471_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2471_In1_c19,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_copy2472_c19);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2471_Out0_copy2472_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In0_c19 <= "" & bh2012_wm2_0_c19 & bh2012_wm2_1_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c0 <= "" & bh2012_wm1_0_c0;
   bh2012_wm2_3_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_c19(0);
   bh2012_wm1_1_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_c19(1);
   Compressor_14_3_Freq300_uid2288_uid2473: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2473_In1_c19,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_copy2474_c19);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2473_Out0_copy2474_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2475_In0_c22 <= "" & bh2012_wm48_4_c22 & bh2012_wm48_5_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2475_In1_c22 <= "" & bh2012_wm47_3_c22;
   bh2012_wm48_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_c22(0);
   bh2012_wm47_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_c22(1);
   bh2012_wm46_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2475: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2475_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2475_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_copy2476_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2475_Out0_copy2476_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2477_In0_c22 <= "" & bh2012_wm46_4_c22 & bh2012_wm46_5_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2477_In1_c22 <= "" & bh2012_wm45_5_c22;
   bh2012_wm46_7_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_c22(0);
   bh2012_wm45_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_c22(1);
   bh2012_wm44_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2477: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2477_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2477_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_copy2478_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2477_Out0_copy2478_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2479_In0_c22 <= "" & bh2012_wm44_4_c22 & bh2012_wm44_5_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2479_In1_c22 <= "" & bh2012_wm43_6_c22 & bh2012_wm43_7_c22;
   bh2012_wm44_7_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_c22(0);
   bh2012_wm43_8_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_c22(1);
   bh2012_wm42_9_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2479: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2479_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2479_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_copy2480_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2479_Out0_copy2480_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2481_In0_c22 <= "" & bh2012_wm41_9_c22 & bh2012_wm41_10_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2481_In1_c22 <= "" & bh2012_wm40_10_c22 & bh2012_wm40_11_c22;
   bh2012_wm41_11_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_c22(0);
   bh2012_wm40_12_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_c22(1);
   bh2012_wm39_15_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2481: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2481_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2481_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_copy2482_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2481_Out0_copy2482_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2483_In0_c22 <= "" & bh2012_wm39_13_c22 & bh2012_wm39_14_c22 & "0";
   bh2012_wm39_16_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_c22(0);
   bh2012_wm38_16_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_c22(1);
   Compressor_3_2_Freq300_uid2264_uid2483: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2483_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_copy2484_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_c22 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2483_Out0_copy2484_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2485_In0_c22 <= "" & bh2012_wm38_12_c22 & bh2012_wm38_13_c22 & bh2012_wm38_14_c22 & bh2012_wm38_15_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2485_In1_c22 <= "" & bh2012_wm37_15_c22;
   bh2012_wm38_17_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_c22(0);
   bh2012_wm37_17_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_c22(1);
   bh2012_wm36_19_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2485: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2485_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2485_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_copy2486_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2485_Out0_copy2486_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In0_c22 <= "" & bh2012_wm36_15_c22 & bh2012_wm36_16_c22 & bh2012_wm36_17_c22 & bh2012_wm36_18_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c0 <= "" & "0";
   bh2012_wm36_20_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_c22(0);
   bh2012_wm35_20_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_c22(1);
   bh2012_wm34_18_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2487: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2487_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_copy2488_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2487_Out0_copy2488_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2489_In0_c22 <= "" & bh2012_wm35_17_c22 & bh2012_wm35_18_c22 & bh2012_wm35_19_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2489_In1_c22 <= "" & bh2012_wm34_16_c22 & bh2012_wm34_17_c22;
   bh2012_wm35_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_c23(0);
   bh2012_wm34_19_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_c23(1);
   bh2012_wm33_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2489: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2489_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2489_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_copy2490_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2489_Out0_copy2490_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In0_c22 <= "" & bh2012_wm33_18_c22 & bh2012_wm33_19_c22 & bh2012_wm33_20_c22 & bh2012_wm33_21_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c0 <= "" & "0";
   bh2012_wm33_23_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_c23(0);
   bh2012_wm32_20_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_c23(1);
   bh2012_wm31_20_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2491: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2491_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_copy2492_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2491_Out0_copy2492_c23; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2493_In0_c22 <= "" & bh2012_wm32_17_c22 & bh2012_wm32_18_c22 & bh2012_wm32_19_c22;
   bh2012_wm32_21_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_c23(0);
   bh2012_wm31_21_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_c23(1);
   Compressor_3_2_Freq300_uid2264_uid2493: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2493_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_copy2494_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2493_Out0_copy2494_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2495_In0_c22 <= "" & bh2012_wm31_17_c22 & bh2012_wm31_18_c22 & bh2012_wm31_19_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2495_In1_c22 <= "" & bh2012_wm30_18_c22 & bh2012_wm30_19_c22;
   bh2012_wm31_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_c23(0);
   bh2012_wm30_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_c23(1);
   bh2012_wm29_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2495: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2495_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2495_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_copy2496_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2495_Out0_copy2496_c23; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2497_In0_c22 <= "" & bh2012_wm29_18_c22 & bh2012_wm29_19_c22 & bh2012_wm29_20_c22;
   bh2012_wm29_22_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_c23(0);
   bh2012_wm28_20_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_c23(1);
   Compressor_3_2_Freq300_uid2264_uid2497: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2497_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_copy2498_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2497_Out0_copy2498_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In0_c22 <= "" & bh2012_wm28_16_c22 & bh2012_wm28_17_c22 & bh2012_wm28_18_c22 & bh2012_wm28_19_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c0 <= "" & "0";
   bh2012_wm28_21_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_c23(0);
   bh2012_wm27_20_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_c23(1);
   bh2012_wm26_20_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2499: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2499_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_copy2500_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2499_Out0_copy2500_c23; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2501_In0_c22 <= "" & bh2012_wm27_17_c22 & bh2012_wm27_18_c22 & bh2012_wm27_19_c22;
   bh2012_wm27_21_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_c23(0);
   bh2012_wm26_21_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_c23(1);
   Compressor_3_2_Freq300_uid2264_uid2501: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2501_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_copy2502_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2501_Out0_copy2502_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2503_In0_c22 <= "" & bh2012_wm26_17_c22 & bh2012_wm26_18_c22 & bh2012_wm26_19_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2503_In1_c22 <= "" & bh2012_wm25_17_c22 & bh2012_wm25_18_c22;
   bh2012_wm26_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_c23(0);
   bh2012_wm25_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_c23(1);
   bh2012_wm24_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2503: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2503_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2503_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_copy2504_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2503_Out0_copy2504_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2505_In0_c22 <= "" & bh2012_wm24_17_c22 & bh2012_wm24_18_c22 & bh2012_wm24_19_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2505_In1_c22 <= "" & bh2012_wm23_17_c22 & bh2012_wm23_18_c22;
   bh2012_wm24_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_c23(0);
   bh2012_wm23_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_c23(1);
   bh2012_wm22_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2505: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2505_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2505_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_copy2506_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2505_Out0_copy2506_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In0_c22 <= "" & bh2012_wm22_16_c22 & bh2012_wm22_17_c22 & bh2012_wm22_18_c22 & bh2012_wm22_19_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c0 <= "" & "0";
   bh2012_wm22_21_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_c22(0);
   bh2012_wm21_21_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_c22(1);
   bh2012_wm20_17_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2507: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2507_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_copy2508_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2507_Out0_copy2508_c22; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2509_In0_c22 <= "" & bh2012_wm21_18_c22 & bh2012_wm21_19_c22 & bh2012_wm21_20_c22;
   bh2012_wm21_22_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_c23(0);
   bh2012_wm20_18_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_c23(1);
   Compressor_3_2_Freq300_uid2264_uid2509: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2509_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_copy2510_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2509_Out0_copy2510_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In0_c22 <= "" & bh2012_wm20_13_c22 & bh2012_wm20_14_c22 & bh2012_wm20_15_c22 & bh2012_wm20_16_c22;
   Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c0 <= "" & "0";
   bh2012_wm20_19_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_c23(0);
   bh2012_wm19_20_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_c23(1);
   bh2012_wm18_19_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2511: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2511_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_copy2512_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2511_Out0_copy2512_c23; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2513_In0_c22 <= "" & bh2012_wm19_17_c22 & bh2012_wm19_18_c22 & bh2012_wm19_19_c22;
   bh2012_wm19_21_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_c23(0);
   bh2012_wm18_20_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_c23(1);
   Compressor_3_2_Freq300_uid2264_uid2513: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2513_In0_c22,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_copy2514_c22);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2513_Out0_copy2514_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2515_In0_c22 <= "" & bh2012_wm18_16_c22 & bh2012_wm18_17_c22 & bh2012_wm18_18_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2515_In1_c22 <= "" & bh2012_wm17_15_c22 & bh2012_wm17_16_c22;
   bh2012_wm18_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_c23(0);
   bh2012_wm17_18_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_c23(1);
   bh2012_wm16_18_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2515: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2515_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2515_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_copy2516_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2515_Out0_copy2516_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2517_In0_c22 <= "" & bh2012_wm16_15_c22 & bh2012_wm16_16_c22 & bh2012_wm16_17_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2517_In1_c22 <= "" & bh2012_wm15_12_c22 & bh2012_wm15_13_c22;
   bh2012_wm16_19_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_c23(0);
   bh2012_wm15_15_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_c23(1);
   bh2012_wm14_14_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2517: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2517_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2517_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_copy2518_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2517_Out0_copy2518_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2519_In0_c22 <= "" & bh2012_wm14_11_c22 & bh2012_wm14_12_c22 & bh2012_wm14_13_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2519_In1_c22 <= "" & bh2012_wm13_9_c22 & bh2012_wm13_10_c22;
   bh2012_wm14_15_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_c23(0);
   bh2012_wm13_12_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_c23(1);
   bh2012_wm12_12_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2519: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2519_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2519_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_copy2520_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2519_Out0_copy2520_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2521_In0_c22 <= "" & bh2012_wm12_9_c22 & bh2012_wm12_10_c22 & bh2012_wm12_11_c22;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2521_In1_c22 <= "" & bh2012_wm11_6_c22 & bh2012_wm11_7_c22;
   bh2012_wm12_13_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_c22(0);
   bh2012_wm11_8_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_c22(1);
   bh2012_wm10_9_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2521: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2521_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2521_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_copy2522_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2521_Out0_copy2522_c22; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2523_In0_c22 <= "" & bh2012_wm10_7_c22 & bh2012_wm10_8_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2523_In1_c22 <= "" & bh2012_wm9_4_c22 & bh2012_wm9_5_c22;
   bh2012_wm10_10_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_c22(0);
   bh2012_wm9_6_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_c22(1);
   bh2012_wm8_6_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_c22(2);
   Compressor_23_3_Freq300_uid2256_uid2523: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2523_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2523_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_copy2524_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_c22 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2523_Out0_copy2524_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2525_In0_c22 <= "" & bh2012_wm8_4_c22 & bh2012_wm8_5_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2525_In1_c22 <= "" & bh2012_wm7_3_c22;
   bh2012_wm8_7_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_c22(0);
   bh2012_wm7_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_c22(1);
   bh2012_wm6_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2525: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2525_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2525_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_copy2526_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2525_Out0_copy2526_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2527_In0_c22 <= "" & bh2012_wm6_4_c22 & bh2012_wm6_5_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2527_In1_c22 <= "" & bh2012_wm5_3_c22;
   bh2012_wm6_7_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_c22(0);
   bh2012_wm5_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_c22(1);
   bh2012_wm4_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2527: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2527_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2527_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_copy2528_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2527_Out0_copy2528_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In0_c22 <= "" & bh2012_wm4_4_c22 & bh2012_wm4_5_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c19 <= "" & bh2012_wm3_3_c19;
   bh2012_wm4_7_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_c22(0);
   bh2012_wm3_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_c22(1);
   bh2012_wm2_4_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2529: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2529_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_copy2530_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2529_Out0_copy2530_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2531_In0_c19 <= "" & bh2012_wm2_2_c19 & bh2012_wm2_3_c19 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2531_In1_c19 <= "" & bh2012_wm1_1_c19;
   bh2012_wm2_5_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_c19(0);
   bh2012_wm1_2_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_c19(1);
   Compressor_14_3_Freq300_uid2288_uid2531: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2531_In0_c19,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2531_In1_c19,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_copy2532_c19);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_c19 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2531_Out0_copy2532_c19; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2533_In0_c22 <= "" & bh2012_wm46_6_c22 & bh2012_wm46_7_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2533_In1_c22 <= "" & bh2012_wm45_6_c22;
   bh2012_wm46_8_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_c23(0);
   bh2012_wm45_7_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_c23(1);
   bh2012_wm44_8_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2533: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2533_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2533_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_copy2534_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2533_Out0_copy2534_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2535_In0_c22 <= "" & bh2012_wm44_6_c22 & bh2012_wm44_7_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2535_In1_c22 <= "" & bh2012_wm43_8_c22;
   bh2012_wm44_9_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_c23(0);
   bh2012_wm43_9_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_c23(1);
   bh2012_wm42_10_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2535: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2535_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2535_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_copy2536_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2535_Out0_copy2536_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2537_In0_c22 <= "" & bh2012_wm42_8_c22 & bh2012_wm42_9_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2537_In1_c22 <= "" & bh2012_wm41_11_c22;
   bh2012_wm42_11_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_c23(0);
   bh2012_wm41_12_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_c23(1);
   bh2012_wm40_13_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2537: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2537_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2537_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_copy2538_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2537_Out0_copy2538_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2539_In0_c22 <= "" & bh2012_wm39_15_c22 & bh2012_wm39_16_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2539_In1_c22 <= "" & bh2012_wm38_16_c22 & bh2012_wm38_17_c22;
   bh2012_wm39_17_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_c23(0);
   bh2012_wm38_18_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_c23(1);
   bh2012_wm37_18_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2539: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2539_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2539_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_copy2540_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2539_Out0_copy2540_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2541_In0_c22 <= "" & bh2012_wm37_16_c22 & bh2012_wm37_17_c22 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2541_In1_c22 <= "" & bh2012_wm36_19_c22 & bh2012_wm36_20_c22;
   bh2012_wm37_19_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_c23(0);
   bh2012_wm36_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_c23(1);
   bh2012_wm35_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2541: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2541_In0_c22,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2541_In1_c22,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_copy2542_c22);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2541_Out0_copy2542_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2543_In0_c23 <= "" & bh2012_wm35_20_c23 & bh2012_wm35_21_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2543_In1_c23 <= "" & bh2012_wm34_18_c23 & bh2012_wm34_19_c23;
   bh2012_wm35_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_c23(0);
   bh2012_wm34_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_c23(1);
   bh2012_wm33_24_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2543: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2543_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2543_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_copy2544_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2543_Out0_copy2544_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2545_In0_c23 <= "" & bh2012_wm33_22_c23 & bh2012_wm33_23_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2545_In1_c23 <= "" & bh2012_wm32_20_c23 & bh2012_wm32_21_c23;
   bh2012_wm33_25_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_c23(0);
   bh2012_wm32_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_c23(1);
   bh2012_wm31_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2545: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2545_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2545_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_copy2546_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2545_Out0_copy2546_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2547_In0_c23 <= "" & bh2012_wm31_20_c23 & bh2012_wm31_21_c23 & bh2012_wm31_22_c23;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2547_In1_c23 <= "" & bh2012_wm30_20_c23 & bh2012_wm30_21_c23;
   bh2012_wm31_24_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_c23(0);
   bh2012_wm30_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_c23(1);
   bh2012_wm29_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2547: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2547_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2547_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_copy2548_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2547_Out0_copy2548_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2549_In0_c23 <= "" & bh2012_wm29_21_c23 & bh2012_wm29_22_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2549_In1_c23 <= "" & bh2012_wm28_20_c23 & bh2012_wm28_21_c23;
   bh2012_wm29_24_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_c23(0);
   bh2012_wm28_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_c23(1);
   bh2012_wm27_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2549: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2549_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2549_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_copy2550_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2549_Out0_copy2550_c23; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2264_bh2012_uid2551_In0_c23 <= "" & bh2012_wm27_20_c23 & bh2012_wm27_21_c23 & "0";
   bh2012_wm27_23_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_c23(0);
   bh2012_wm26_23_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_c23(1);
   Compressor_3_2_Freq300_uid2264_uid2551: Compressor_3_2_Freq300_uid2264
      port map ( X0 => Compressor_3_2_Freq300_uid2264_bh2012_uid2551_In0_c23,
                 R => Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_copy2552_c23);
   Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_c23 <= Compressor_3_2_Freq300_uid2264_bh2012_uid2551_Out0_copy2552_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2553_In0_c23 <= "" & bh2012_wm26_20_c23 & bh2012_wm26_21_c23 & bh2012_wm26_22_c23;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2553_In1_c23 <= "" & bh2012_wm25_19_c23 & bh2012_wm25_20_c23;
   bh2012_wm26_24_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_c23(0);
   bh2012_wm25_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_c23(1);
   bh2012_wm24_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2553: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2553_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2553_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_copy2554_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2553_Out0_copy2554_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2555_In0_c23 <= "" & bh2012_wm24_20_c23 & bh2012_wm24_21_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2555_In1_c23 <= "" & bh2012_wm23_19_c23 & bh2012_wm23_20_c23;
   bh2012_wm24_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_c23(0);
   bh2012_wm23_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_c23(1);
   bh2012_wm22_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2555: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2555_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2555_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_copy2556_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2555_Out0_copy2556_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2557_In0_c23 <= "" & bh2012_wm22_20_c23 & bh2012_wm22_21_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2557_In1_c23 <= "" & bh2012_wm21_21_c23 & bh2012_wm21_22_c23;
   bh2012_wm22_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_c23(0);
   bh2012_wm21_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_c23(1);
   bh2012_wm20_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2557: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2557_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2557_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_copy2558_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2557_Out0_copy2558_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2559_In0_c23 <= "" & bh2012_wm20_17_c23 & bh2012_wm20_18_c23 & bh2012_wm20_19_c23;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2559_In1_c23 <= "" & bh2012_wm19_20_c23 & bh2012_wm19_21_c23;
   bh2012_wm20_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_c23(0);
   bh2012_wm19_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_c23(1);
   bh2012_wm18_22_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2559: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2559_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2559_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_copy2560_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2559_Out0_copy2560_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2561_In0_c23 <= "" & bh2012_wm18_19_c23 & bh2012_wm18_20_c23 & bh2012_wm18_21_c23;
   Compressor_23_3_Freq300_uid2256_bh2012_uid2561_In1_c23 <= "" & bh2012_wm17_17_c23 & bh2012_wm17_18_c23;
   bh2012_wm18_23_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_c23(0);
   bh2012_wm17_19_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_c23(1);
   bh2012_wm16_20_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2561: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2561_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2561_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_copy2562_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2561_Out0_copy2562_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2563_In0_c23 <= "" & bh2012_wm16_18_c23 & bh2012_wm16_19_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2563_In1_c23 <= "" & bh2012_wm15_14_c23 & bh2012_wm15_15_c23;
   bh2012_wm16_21_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_c23(0);
   bh2012_wm15_16_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_c23(1);
   bh2012_wm14_16_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2563: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2563_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2563_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_copy2564_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2563_Out0_copy2564_c23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2256_bh2012_uid2565_In0_c23 <= "" & bh2012_wm14_14_c23 & bh2012_wm14_15_c23 & "0";
   Compressor_23_3_Freq300_uid2256_bh2012_uid2565_In1_c23 <= "" & bh2012_wm13_11_c23 & bh2012_wm13_12_c23;
   bh2012_wm14_17_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_c23(0);
   bh2012_wm13_13_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_c23(1);
   bh2012_wm12_14_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_c23(2);
   Compressor_23_3_Freq300_uid2256_uid2565: Compressor_23_3_Freq300_uid2256
      port map ( X0 => Compressor_23_3_Freq300_uid2256_bh2012_uid2565_In0_c23,
                 X1 => Compressor_23_3_Freq300_uid2256_bh2012_uid2565_In1_c23,
                 R => Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_copy2566_c23);
   Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_c23 <= Compressor_23_3_Freq300_uid2256_bh2012_uid2565_Out0_copy2566_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In0_c23 <= "" & bh2012_wm12_12_c23 & bh2012_wm12_13_c23 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In1_c22 <= "" & bh2012_wm11_8_c22;
   bh2012_wm12_15_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_c23(0);
   bh2012_wm11_9_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_c23(1);
   bh2012_wm10_11_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_c23(2);
   Compressor_14_3_Freq300_uid2288_uid2567: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In0_c23,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2567_In1_c23,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_copy2568_c23);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_c23 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2567_Out0_copy2568_c23; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2569_In0_c22 <= "" & bh2012_wm10_9_c22 & bh2012_wm10_10_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2569_In1_c22 <= "" & bh2012_wm9_6_c22;
   bh2012_wm10_12_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_c22(0);
   bh2012_wm9_7_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_c22(1);
   bh2012_wm8_8_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2569: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2569_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2569_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_copy2570_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2569_Out0_copy2570_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2571_In0_c22 <= "" & bh2012_wm8_6_c22 & bh2012_wm8_7_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2571_In1_c22 <= "" & bh2012_wm7_4_c22;
   bh2012_wm8_9_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_c22(0);
   bh2012_wm7_5_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_c22(1);
   bh2012_wm6_8_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2571: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2571_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2571_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_copy2572_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2571_Out0_copy2572_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2573_In0_c22 <= "" & bh2012_wm6_6_c22 & bh2012_wm6_7_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2573_In1_c22 <= "" & bh2012_wm5_4_c22;
   bh2012_wm6_9_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_c22(0);
   bh2012_wm5_5_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_c22(1);
   bh2012_wm4_8_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2573: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2573_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2573_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_copy2574_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2573_Out0_copy2574_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2575_In0_c22 <= "" & bh2012_wm4_6_c22 & bh2012_wm4_7_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2575_In1_c22 <= "" & bh2012_wm3_4_c22;
   bh2012_wm4_9_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_c22(0);
   bh2012_wm3_5_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_c22(1);
   bh2012_wm2_6_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_c22(2);
   Compressor_14_3_Freq300_uid2288_uid2575: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2575_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2575_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_copy2576_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2575_Out0_copy2576_c22; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In0_c22 <= "" & bh2012_wm2_4_c22 & bh2012_wm2_5_c22 & "0" & "0";
   Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c19 <= "" & bh2012_wm1_2_c19;
   bh2012_wm2_7_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_c22(0);
   bh2012_wm1_3_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_c22(1);
   Compressor_14_3_Freq300_uid2288_uid2577: Compressor_14_3_Freq300_uid2288
      port map ( X0 => Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In0_c22,
                 X1 => Compressor_14_3_Freq300_uid2288_bh2012_uid2577_In1_c22,
                 R => Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_copy2578_c22);
   Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_c22 <= Compressor_14_3_Freq300_uid2288_bh2012_uid2577_Out0_copy2578_c22; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh2012_24_c23 <= bh2012_wm45_7_c23 & bh2012_wm46_8_c23 & bh2012_wm47_4_c23 & bh2012_wm48_6_c23 & bh2012_wm49_3_c23 & bh2012_wm50_4_c23 & bh2012_wm51_2_c23 & bh2012_wm52_2_c23 & bh2012_wm53_0_c23 & bh2012_wm54_0_c23 & bh2012_wm55_0_c23 & bh2012_wm56_0_c23 & bh2012_wm57_0_c23 & bh2012_wm58_0_c23 & bh2012_wm59_0_c23 & bh2012_wm60_0_c23 & bh2012_wm61_0_c23 & bh2012_wm62_0_c23 & bh2012_wm63_0_c23 & bh2012_wm64_0_c23 & bh2012_wm65_0_c23 & bh2012_wm66_0_c23 & bh2012_wm67_0_c23 & bh2012_wm68_0_c23 & bh2012_wm69_0_c23;

   bitheapFinalAdd_bh2012_In0_c23 <= "0" & bh2012_wm1_3_c23 & bh2012_wm2_6_c23 & bh2012_wm3_5_c23 & bh2012_wm4_8_c23 & bh2012_wm5_5_c23 & bh2012_wm6_8_c23 & bh2012_wm7_5_c23 & bh2012_wm8_8_c23 & bh2012_wm9_7_c23 & bh2012_wm10_11_c23 & bh2012_wm11_9_c23 & bh2012_wm12_14_c23 & bh2012_wm13_13_c23 & bh2012_wm14_16_c23 & bh2012_wm15_16_c23 & bh2012_wm16_20_c23 & bh2012_wm17_19_c23 & bh2012_wm18_22_c23 & bh2012_wm19_22_c23 & bh2012_wm20_20_c23 & bh2012_wm21_23_c23 & bh2012_wm22_22_c23 & bh2012_wm23_21_c23 & bh2012_wm24_22_c23 & bh2012_wm25_21_c23 & bh2012_wm26_23_c23 & bh2012_wm27_22_c23 & bh2012_wm28_22_c23 & bh2012_wm29_23_c23 & bh2012_wm30_22_c23 & bh2012_wm31_23_c23 & bh2012_wm32_22_c23 & bh2012_wm33_24_c23 & bh2012_wm34_20_c23 & bh2012_wm35_22_c23 & bh2012_wm36_21_c23 & bh2012_wm37_18_c23 & bh2012_wm38_18_c23 & bh2012_wm39_17_c23 & bh2012_wm40_12_c23 & bh2012_wm41_12_c23 & bh2012_wm42_10_c23 & bh2012_wm43_9_c23 & bh2012_wm44_8_c23;
   bitheapFinalAdd_bh2012_In1_c23 <= "0" & "0" & bh2012_wm2_7_c23 & "0" & bh2012_wm4_9_c23 & "0" & bh2012_wm6_9_c23 & "0" & bh2012_wm8_9_c23 & "0" & bh2012_wm10_12_c23 & "0" & bh2012_wm12_15_c23 & "0" & bh2012_wm14_17_c23 & "0" & bh2012_wm16_21_c23 & "0" & bh2012_wm18_23_c23 & "0" & bh2012_wm20_21_c23 & "0" & bh2012_wm22_23_c23 & "0" & bh2012_wm24_23_c23 & "0" & bh2012_wm26_24_c23 & bh2012_wm27_23_c23 & "0" & bh2012_wm29_24_c23 & "0" & bh2012_wm31_24_c23 & "0" & bh2012_wm33_25_c23 & "0" & bh2012_wm35_23_c23 & "0" & bh2012_wm37_19_c23 & "0" & "0" & bh2012_wm40_13_c23 & "0" & bh2012_wm42_11_c23 & "0" & bh2012_wm44_9_c23;
   bitheapFinalAdd_bh2012_Cin_c0 <= '0';

   bitheapFinalAdd_bh2012: IntAdder_45_Freq300_uid2580
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 Cin => bitheapFinalAdd_bh2012_Cin_c0,
                 X => bitheapFinalAdd_bh2012_In0_c23,
                 Y => bitheapFinalAdd_bh2012_In1_c23,
                 R => bitheapFinalAdd_bh2012_Out_c23);
   bitheapResult_bh2012_c23 <= bitheapFinalAdd_bh2012_Out_c23(43 downto 0) & tmp_bitheapResult_bh2012_24_c23;
   RR_c23 <= signed(bitheapResult_bh2012_c23(68 downto 28));
R <= std_logic_vector(RR_c23);  
end architecture;

--------------------------------------------------------------------------------
--                     FixHornerEvaluator_Freq300_uid1539
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin (2014-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: Y A0 A1 A2
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixHornerEvaluator_Freq300_uid1539 is
    port (clk, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          Y : in  std_logic_vector(28 downto 0);
          A0 : in  std_logic_vector(39 downto 0);
          A1 : in  std_logic_vector(32 downto 0);
          A2 : in  std_logic_vector(24 downto 0);
          R : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of FixHornerEvaluator_Freq300_uid1539 is
   component FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid1541 is
      port ( clk, ce_20, ce_21 : in std_logic;
             X : in  std_logic_vector(24 downto 0);
             Y : in  std_logic_vector(24 downto 0);
             A : in  std_logic_vector(32 downto 0);
             R : out  std_logic_vector(32 downto 0)   );
   end component;

   component FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid2011 is
      port ( clk, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             X : in  std_logic_vector(28 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             A : in  std_logic_vector(39 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

signal Ys_c19 :  signed(0+28 downto 0);
signal As0_c19 :  signed(-2+41 downto 0);
signal As1_c19 :  signed(-9+41 downto 0);
signal As2_c19 :  signed(-17+41 downto 0);
signal S2_c19 :  signed(-17+41 downto 0);
signal YsTrunc1_c19 :  signed(0+24 downto 0);
signal SS1_c21 :  std_logic_vector(32 downto 0);
signal S1_c21 :  signed(-9+41 downto 0);
signal YsTrunc0_c19 :  signed(0+28 downto 0);
signal SS0_c23 :  std_logic_vector(40 downto 0);
signal S0_c23 :  signed(-1+41 downto 0);
signal Rs_c23 :  signed(-2+37 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
            end if;
            if ce_21 = '1' then
            end if;
            if ce_22 = '1' then
            end if;
            if ce_23 = '1' then
            end if;
         end if;
      end process;
   Ys_c19 <= signed(Y);
   As0_c19 <= signed(A0);
   As1_c19 <= signed(A1);
   As2_c19 <= signed(A2);
   S2_c19 <= As2_c19(24 downto 0); -- fix resize from (-17, -41) to (-17, -41)
   YsTrunc1_c19 <= Ys_c19(28 downto 4); -- fix resize from (0, -28) to (0, -24)
   FixHornerEvaluator_Freq300_uid1539_step_1: FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid1541
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 A => std_logic_vector(As1_c19),
                 X => std_logic_vector(YsTrunc1_c19),
                 Y => std_logic_vector(S2_c19),
                 R => SS1_c21);
S1_c21 <= signed(SS1_c21);
   YsTrunc0_c19 <= Ys_c19(28 downto 0); -- fix resize from (0, -28) to (0, -28)
   FixHornerEvaluator_Freq300_uid1539_step_0: FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid2011
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 A => std_logic_vector(As0_c19),
                 X => std_logic_vector(YsTrunc0_c19),
                 Y => std_logic_vector(S1_c21),
                 R => SS0_c23);
S0_c23 <= signed(SS0_c23);
   Rs_c23 <= S0_c23(39 downto 4); -- fix resize from (-1, -41) to (-2, -37)
   R <= std_logic_vector(Rs_c23);
end architecture;

--------------------------------------------------------------------------------
--                 FixFunctionByPiecewisePoly_Freq300_uid1534
-- Evaluator for 1b19*(exp(x*1b-10)-x*1b-10-1) on [0,1) for lsbIn=-36 (wIn=36), msbout=-2, lsbOut=-37 (wOut=36). Out interval: [0; 0.250081]. Output is unsigned

-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2014-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByPiecewisePoly_Freq300_uid1534 is
    port (clk, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          X : in  std_logic_vector(35 downto 0);
          Y : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of FixFunctionByPiecewisePoly_Freq300_uid1534 is
   component coeffTable_Freq300_uid1536 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(94 downto 0)   );
   end component;

   component FixHornerEvaluator_Freq300_uid1539 is
      port ( clk, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             Y : in  std_logic_vector(28 downto 0);
             A0 : in  std_logic_vector(39 downto 0);
             A1 : in  std_logic_vector(32 downto 0);
             A2 : in  std_logic_vector(24 downto 0);
             R : out  std_logic_vector(35 downto 0)   );
   end component;

signal A_c19 :  std_logic_vector(6 downto 0);
signal Z_c19 :  std_logic_vector(28 downto 0);
signal Zs_c19 :  std_logic_vector(28 downto 0);
signal Coeffs_c19 :  std_logic_vector(94 downto 0);
signal Coeffs_copy1537_c19 :  std_logic_vector(94 downto 0);
signal A2_c19 :  std_logic_vector(24 downto 0);
signal A1_c19 :  std_logic_vector(32 downto 0);
signal A0_c19 :  std_logic_vector(39 downto 0);
signal HornerOutput_c23 :  std_logic_vector(35 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_20 = '1' then
            end if;
            if ce_21 = '1' then
            end if;
            if ce_22 = '1' then
            end if;
            if ce_23 = '1' then
            end if;
         end if;
      end process;
   A_c19 <= X(35 downto 29);
   Z_c19 <= X(28 downto 0);
   Zs_c19 <= (not Z_c19(28)) & Z_c19(27 downto 0); -- centering the interval
   coeffTable: coeffTable_Freq300_uid1536
      port map ( X => A_c19,
                 Y => Coeffs_copy1537_c19);
   Coeffs_c19 <= Coeffs_copy1537_c19; -- output copy to hold a pipeline register if needed
   --  Split the table output into each coefficient, adding back the constant signs if any
   A2_c19 <= "0" & Coeffs_c19(23 downto 0);
   A1_c19 <= "0" & Coeffs_c19(55 downto 24);
   A0_c19 <= "0" & Coeffs_c19(94 downto 56);
   Horner: FixHornerEvaluator_Freq300_uid1539
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 A0 => A0_c19,
                 A1 => A1_c19,
                 A2 => A2_c19,
                 Y => Zs_c19,
                 R => HornerOutput_c23);
   Y <= std_logic_vector(HornerOutput_c23);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_47_Freq300_uid2583
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_47_Freq300_uid2583 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(46 downto 0);
          Y : in  std_logic_vector(46 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(46 downto 0)   );
end entity;

architecture arch of IntAdder_47_Freq300_uid2583 is
signal Rtmp_c24 :  std_logic_vector(46 downto 0);
signal X_c20, X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(46 downto 0);
signal Y_c24 :  std_logic_vector(46 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19, Cin_c20, Cin_c21, Cin_c22, Cin_c23, Cin_c24 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               Cin_c19 <= Cin_c18;
            end if;
            if ce_20 = '1' then
               X_c20 <= X;
               Cin_c20 <= Cin_c19;
            end if;
            if ce_21 = '1' then
               X_c21 <= X_c20;
               Cin_c21 <= Cin_c20;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
               Cin_c22 <= Cin_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
               Cin_c23 <= Cin_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
               Y_c24 <= Y;
               Cin_c24 <= Cin_c23;
            end if;
         end if;
      end process;
   Rtmp_c24 <= X_c24 + Y_c24 + Cin_c24;
   R <= Rtmp_c24;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid2589
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid2589 is
    port (clk, ce_21, ce_22, ce_23, ce_24, ce_25 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid2589 is
signal Mfull_c24, Mfull_c25 :  std_logic_vector(40 downto 0);
signal M_c25 :  std_logic_vector(40 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
            if ce_25 = '1' then
               Mfull_c25 <= Mfull_c24;
            end if;
         end if;
      end process;
   Mfull_c24 <= std_logic_vector(unsigned(X_c24) * unsigned(Y)); -- multiplier
   M_c25 <= Mfull_c25(40 downto 0);
   R <= M_c25;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2591
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2591 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2591 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2593
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2593 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2593 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2595
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2595 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2595 is
   component MultTable_Freq300_uid2597 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(3 downto 0);
signal Y1_c24 :  std_logic_vector(3 downto 0);
signal Y1_copy2598_c24 :  std_logic_vector(3 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2597
      port map ( X => Xtable_c24,
                 Y => Y1_copy2598_c24);
   Y1_c24 <= Y1_copy2598_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2600
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2600 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2600 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid2602
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid2602 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid2602 is
signal replicated_c24 :  std_logic_vector(1 downto 0);
signal prod_c24 :  std_logic_vector(1 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
   replicated_c24 <= (1 downto 0 => Y(0));
   prod_c24 <= X_c24 and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2604
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2604 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2604 is
   component MultTable_Freq300_uid2606 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2607_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2606
      port map ( X => Xtable_c24,
                 Y => Y1_copy2607_c24);
   Y1_c24 <= Y1_copy2607_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2609
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2609 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2609 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2611
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2611 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2611 is
   component MultTable_Freq300_uid2613 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2614_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2613
      port map ( X => Xtable_c24,
                 Y => Y1_copy2614_c24);
   Y1_c24 <= Y1_copy2614_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2616
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2616 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2616 is
   component MultTable_Freq300_uid2618 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2619_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2618
      port map ( X => Xtable_c24,
                 Y => Y1_copy2619_c24);
   Y1_c24 <= Y1_copy2619_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2621
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2621 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2621 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2623
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2623 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2623 is
   component MultTable_Freq300_uid2625 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(3 downto 0);
signal Y1_c24 :  std_logic_vector(3 downto 0);
signal Y1_copy2626_c24 :  std_logic_vector(3 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2625
      port map ( X => Xtable_c24,
                 Y => Y1_copy2626_c24);
   Y1_c24 <= Y1_copy2626_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2628
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2628 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2628 is
   component MultTable_Freq300_uid2630 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2631_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2630
      port map ( X => Xtable_c24,
                 Y => Y1_copy2631_c24);
   Y1_c24 <= Y1_copy2631_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2633
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2633 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2633 is
   component MultTable_Freq300_uid2635 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2636_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2635
      port map ( X => Xtable_c24,
                 Y => Y1_copy2636_c24);
   Y1_c24 <= Y1_copy2636_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2638
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2638 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2638 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid2640
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid2640 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid2640 is
signal replicated_c24 :  std_logic_vector(1 downto 0);
signal prod_c24 :  std_logic_vector(1 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
   replicated_c24 <= (1 downto 0 => Y(0));
   prod_c24 <= X_c24 and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2642
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2642 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2642 is
   component MultTable_Freq300_uid2644 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2645_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2644
      port map ( X => Xtable_c24,
                 Y => Y1_copy2645_c24);
   Y1_c24 <= Y1_copy2645_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2647
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2647 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2647 is
   component MultTable_Freq300_uid2649 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2650_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2649
      port map ( X => Xtable_c24,
                 Y => Y1_copy2650_c24);
   Y1_c24 <= Y1_copy2650_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2652
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2652 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2652 is
   component MultTable_Freq300_uid2654 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2655_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2654
      port map ( X => Xtable_c24,
                 Y => Y1_copy2655_c24);
   Y1_c24 <= Y1_copy2655_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2657
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2657 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2657 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2659
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2659 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2659 is
   component MultTable_Freq300_uid2661 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2662_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2661
      port map ( X => Xtable_c24,
                 Y => Y1_copy2662_c24);
   Y1_c24 <= Y1_copy2662_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2664
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2664 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2664 is
   component MultTable_Freq300_uid2666 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2667_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2666
      port map ( X => Xtable_c24,
                 Y => Y1_copy2667_c24);
   Y1_c24 <= Y1_copy2667_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2669
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2669 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2669 is
   component MultTable_Freq300_uid2671 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2672_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2671
      port map ( X => Xtable_c24,
                 Y => Y1_copy2672_c24);
   Y1_c24 <= Y1_copy2672_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2674
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2674 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2674 is
   component MultTable_Freq300_uid2676 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2677_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2676
      port map ( X => Xtable_c24,
                 Y => Y1_copy2677_c24);
   Y1_c24 <= Y1_copy2677_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x23_Freq300_uid2679
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x23_Freq300_uid2679 is
    port (clk, ce_21, ce_22, ce_23, ce_24, ce_25 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(22 downto 0);
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of DSPBlock_17x23_Freq300_uid2679 is
signal Mfull_c24, Mfull_c25 :  std_logic_vector(39 downto 0);
signal M_c25 :  std_logic_vector(39 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
            if ce_25 = '1' then
               Mfull_c25 <= Mfull_c24;
            end if;
         end if;
      end process;
   Mfull_c24 <= std_logic_vector(unsigned(X_c24) * unsigned(Y)); -- multiplier
   M_c25 <= Mfull_c25(39 downto 0);
   R <= M_c25;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x23_Freq300_uid2681
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x23_Freq300_uid2681 is
    port (clk, ce_21, ce_22, ce_23, ce_24, ce_25 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(22 downto 0);
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of DSPBlock_17x23_Freq300_uid2681 is
signal Mfull_c24, Mfull_c25 :  std_logic_vector(39 downto 0);
signal M_c25 :  std_logic_vector(39 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
            if ce_25 = '1' then
               Mfull_c25 <= Mfull_c24;
            end if;
         end if;
      end process;
   Mfull_c24 <= std_logic_vector(unsigned(X_c24) * unsigned(Y)); -- multiplier
   M_c25 <= Mfull_c25(39 downto 0);
   R <= M_c25;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2683
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2683 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2683 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2685
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2685 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2685 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2687
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2687 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2687 is
   component MultTable_Freq300_uid2689 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(3 downto 0);
signal Y1_c24 :  std_logic_vector(3 downto 0);
signal Y1_copy2690_c24 :  std_logic_vector(3 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2689
      port map ( X => Xtable_c24,
                 Y => Y1_copy2690_c24);
   Y1_c24 <= Y1_copy2690_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2692
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2692 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2692 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid2694
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid2694 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid2694 is
signal replicated_c24 :  std_logic_vector(1 downto 0);
signal prod_c24 :  std_logic_vector(1 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
   replicated_c24 <= (1 downto 0 => Y(0));
   prod_c24 <= X_c24 and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2696
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2696 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2696 is
   component MultTable_Freq300_uid2698 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2699_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2698
      port map ( X => Xtable_c24,
                 Y => Y1_copy2699_c24);
   Y1_c24 <= Y1_copy2699_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2701
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2701 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2701 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2703
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2703 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2703 is
   component MultTable_Freq300_uid2705 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2706_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2705
      port map ( X => Xtable_c24,
                 Y => Y1_copy2706_c24);
   Y1_c24 <= Y1_copy2706_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2708
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2708 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2708 is
   component MultTable_Freq300_uid2710 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2711_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2710
      port map ( X => Xtable_c24,
                 Y => Y1_copy2711_c24);
   Y1_c24 <= Y1_copy2711_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2713
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2713 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2713 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid2715
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid2715 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid2715 is
   component MultTable_Freq300_uid2717 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(3 downto 0);
signal Y1_c24 :  std_logic_vector(3 downto 0);
signal Y1_copy2718_c24 :  std_logic_vector(3 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2717
      port map ( X => Xtable_c24,
                 Y => Y1_copy2718_c24);
   Y1_c24 <= Y1_copy2718_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2720
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2720 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2720 is
   component MultTable_Freq300_uid2722 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2723_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2722
      port map ( X => Xtable_c24,
                 Y => Y1_copy2723_c24);
   Y1_c24 <= Y1_copy2723_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2725
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2725 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2725 is
   component MultTable_Freq300_uid2727 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2728_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2727
      port map ( X => Xtable_c24,
                 Y => Y1_copy2728_c24);
   Y1_c24 <= Y1_copy2728_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid2730
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid2730 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid2730 is
signal replicated_c20, replicated_c21, replicated_c22, replicated_c23, replicated_c24 :  std_logic_vector(0 downto 0);
signal prod_c24 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               replicated_c21 <= replicated_c20;
            end if;
            if ce_22 = '1' then
               replicated_c22 <= replicated_c21;
            end if;
            if ce_23 = '1' then
               replicated_c23 <= replicated_c22;
            end if;
            if ce_24 = '1' then
               replicated_c24 <= replicated_c23;
            end if;
         end if;
      end process;
   replicated_c20 <= (0 downto 0 => X(0));
   prod_c24 <= Y and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid2732
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid2732 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid2732 is
signal replicated_c24 :  std_logic_vector(1 downto 0);
signal prod_c24 :  std_logic_vector(1 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
   replicated_c24 <= (1 downto 0 => Y(0));
   prod_c24 <= X_c24 and replicated_c24;
   R <= prod_c24;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2734
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2734 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2734 is
   component MultTable_Freq300_uid2736 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2737_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2736
      port map ( X => Xtable_c24,
                 Y => Y1_copy2737_c24);
   Y1_c24 <= Y1_copy2737_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2739
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2739 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2739 is
   component MultTable_Freq300_uid2741 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2742_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2741
      port map ( X => Xtable_c24,
                 Y => Y1_copy2742_c24);
   Y1_c24 <= Y1_copy2742_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2744
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2744 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2744 is
   component MultTable_Freq300_uid2746 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2747_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2746
      port map ( X => Xtable_c24,
                 Y => Y1_copy2747_c24);
   Y1_c24 <= Y1_copy2747_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2749
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2749 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2749 is
   component MultTable_Freq300_uid2751 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2752_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2751
      port map ( X => Xtable_c24,
                 Y => Y1_copy2752_c24);
   Y1_c24 <= Y1_copy2752_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2754
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2754 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2754 is
   component MultTable_Freq300_uid2756 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2757_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2756
      port map ( X => Xtable_c24,
                 Y => Y1_copy2757_c24);
   Y1_c24 <= Y1_copy2757_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2759
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2759 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2759 is
   component MultTable_Freq300_uid2761 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2762_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2761
      port map ( X => Xtable_c24,
                 Y => Y1_copy2762_c24);
   Y1_c24 <= Y1_copy2762_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2764
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2764 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2764 is
   component MultTable_Freq300_uid2766 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2767_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2766
      port map ( X => Xtable_c24,
                 Y => Y1_copy2767_c24);
   Y1_c24 <= Y1_copy2767_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2769
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2769 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2769 is
   component MultTable_Freq300_uid2771 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2772_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2771
      port map ( X => Xtable_c24,
                 Y => Y1_copy2772_c24);
   Y1_c24 <= Y1_copy2772_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2774
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2774 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2774 is
   component MultTable_Freq300_uid2776 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2777_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2776
      port map ( X => Xtable_c24,
                 Y => Y1_copy2777_c24);
   Y1_c24 <= Y1_copy2777_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2779
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2779 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2779 is
   component MultTable_Freq300_uid2781 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2782_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2781
      port map ( X => Xtable_c24,
                 Y => Y1_copy2782_c24);
   Y1_c24 <= Y1_copy2782_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2784
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2784 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2784 is
   component MultTable_Freq300_uid2786 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2787_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2786
      port map ( X => Xtable_c24,
                 Y => Y1_copy2787_c24);
   Y1_c24 <= Y1_copy2787_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2789
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2789 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2789 is
   component MultTable_Freq300_uid2791 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2792_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2791
      port map ( X => Xtable_c24,
                 Y => Y1_copy2792_c24);
   Y1_c24 <= Y1_copy2792_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2794
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2794 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2794 is
   component MultTable_Freq300_uid2796 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2797_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2796
      port map ( X => Xtable_c24,
                 Y => Y1_copy2797_c24);
   Y1_c24 <= Y1_copy2797_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2799
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2799 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2799 is
   component MultTable_Freq300_uid2801 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2802_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2801
      port map ( X => Xtable_c24,
                 Y => Y1_copy2802_c24);
   Y1_c24 <= Y1_copy2802_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2804
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2804 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2804 is
   component MultTable_Freq300_uid2806 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2807_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2806
      port map ( X => Xtable_c24,
                 Y => Y1_copy2807_c24);
   Y1_c24 <= Y1_copy2807_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2809
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2809 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2809 is
   component MultTable_Freq300_uid2811 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2812_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2811
      port map ( X => Xtable_c24,
                 Y => Y1_copy2812_c24);
   Y1_c24 <= Y1_copy2812_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2814
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2814 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2814 is
   component MultTable_Freq300_uid2816 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2817_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2816
      port map ( X => Xtable_c24,
                 Y => Y1_copy2817_c24);
   Y1_c24 <= Y1_copy2817_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2819
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2819 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2819 is
   component MultTable_Freq300_uid2821 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2822_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2821
      port map ( X => Xtable_c24,
                 Y => Y1_copy2822_c24);
   Y1_c24 <= Y1_copy2822_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid2824
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid2824 is
    port (clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid2824 is
   component MultTable_Freq300_uid2826 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c24 :  std_logic_vector(4 downto 0);
signal Y1_c24 :  std_logic_vector(4 downto 0);
signal Y1_copy2827_c24 :  std_logic_vector(4 downto 0);
signal X_c21, X_c22, X_c23, X_c24 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               X_c21 <= X;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
            end if;
         end if;
      end process;
Xtable_c24 <= Y & X_c24;
   R <= Y1_c24;
   TableMult: MultTable_Freq300_uid2826
      port map ( X => Xtable_c24,
                 Y => Y1_copy2827_c24);
   Y1_c24 <= Y1_copy2827_c24; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_50_Freq300_uid3174
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_50_Freq300_uid3174 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
          X : in  std_logic_vector(49 downto 0);
          Y : in  std_logic_vector(49 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of IntAdder_50_Freq300_uid3174 is
signal Rtmp_c26 :  std_logic_vector(49 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19, Cin_c20, Cin_c21, Cin_c22, Cin_c23, Cin_c24, Cin_c25, Cin_c26 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               Cin_c19 <= Cin_c18;
            end if;
            if ce_20 = '1' then
               Cin_c20 <= Cin_c19;
            end if;
            if ce_21 = '1' then
               Cin_c21 <= Cin_c20;
            end if;
            if ce_22 = '1' then
               Cin_c22 <= Cin_c21;
            end if;
            if ce_23 = '1' then
               Cin_c23 <= Cin_c22;
            end if;
            if ce_24 = '1' then
               Cin_c24 <= Cin_c23;
            end if;
            if ce_25 = '1' then
               Cin_c25 <= Cin_c24;
            end if;
            if ce_26 = '1' then
               Cin_c26 <= Cin_c25;
            end if;
         end if;
      end process;
   Rtmp_c26 <= X + Y + Cin_c26;
   R <= Rtmp_c26;
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplier_46x47_48_Freq300_uid2585
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_46x47_48_Freq300_uid2585 is
    port (clk, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
          X : in  std_logic_vector(45 downto 0);
          Y : in  std_logic_vector(46 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_46x47_48_Freq300_uid2585 is
   component DSPBlock_17x24_Freq300_uid2589 is
      port ( clk, ce_21, ce_22, ce_23, ce_24, ce_25 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2591 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2593 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2595 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2600 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid2602 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2604 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2609 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2611 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2616 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2621 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2623 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2628 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2633 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2638 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid2640 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2642 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2647 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2652 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2657 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2659 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2664 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2669 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2674 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x23_Freq300_uid2679 is
      port ( clk, ce_21, ce_22, ce_23, ce_24, ce_25 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(22 downto 0);
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component DSPBlock_17x23_Freq300_uid2681 is
      port ( clk, ce_21, ce_22, ce_23, ce_24, ce_25 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(22 downto 0);
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2683 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2685 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2687 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2692 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid2694 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2696 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2701 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2703 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2708 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2713 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid2715 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2720 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2725 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid2730 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid2732 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2734 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2739 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2744 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2749 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2754 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2759 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2764 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2769 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2774 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2779 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2784 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2789 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2794 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2799 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2804 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2809 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2814 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2819 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid2824 is
      port ( clk, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid2830 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid2834 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid2838 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid2848 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid3032 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_50_Freq300_uid3174 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
             X : in  std_logic_vector(49 downto 0);
             Y : in  std_logic_vector(49 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(49 downto 0)   );
   end component;

signal XX_m2586_c20 :  std_logic_vector(45 downto 0);
signal YY_m2586_c24 :  std_logic_vector(46 downto 0);
signal tile_0_X_c20 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c24 :  std_logic_vector(23 downto 0);
signal tile_0_output_c25 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c25 :  unsigned(40-0 downto 0);
signal bh2587_w29_0_c25, bh2587_w29_0_c26 :  std_logic;
signal bh2587_w30_0_c25, bh2587_w30_0_c26 :  std_logic;
signal bh2587_w31_0_c25, bh2587_w31_0_c26 :  std_logic;
signal bh2587_w32_0_c25, bh2587_w32_0_c26 :  std_logic;
signal bh2587_w33_0_c25, bh2587_w33_0_c26 :  std_logic;
signal bh2587_w34_0_c25, bh2587_w34_0_c26 :  std_logic;
signal bh2587_w35_0_c25, bh2587_w35_0_c26 :  std_logic;
signal bh2587_w36_0_c25 :  std_logic;
signal bh2587_w37_0_c25 :  std_logic;
signal bh2587_w38_0_c25 :  std_logic;
signal bh2587_w39_0_c25 :  std_logic;
signal bh2587_w40_0_c25 :  std_logic;
signal bh2587_w41_0_c25 :  std_logic;
signal bh2587_w42_0_c25 :  std_logic;
signal bh2587_w43_0_c25 :  std_logic;
signal bh2587_w44_0_c25 :  std_logic;
signal bh2587_w45_0_c25 :  std_logic;
signal bh2587_w46_0_c25 :  std_logic;
signal bh2587_w47_0_c25 :  std_logic;
signal bh2587_w48_0_c25 :  std_logic;
signal bh2587_w49_0_c25 :  std_logic;
signal bh2587_w50_0_c25 :  std_logic;
signal bh2587_w51_0_c25 :  std_logic;
signal bh2587_w52_0_c25 :  std_logic;
signal bh2587_w53_0_c25 :  std_logic;
signal bh2587_w54_0_c25 :  std_logic;
signal bh2587_w55_0_c25 :  std_logic;
signal bh2587_w56_0_c25 :  std_logic;
signal bh2587_w57_0_c25 :  std_logic;
signal bh2587_w58_0_c25 :  std_logic;
signal bh2587_w59_0_c25 :  std_logic;
signal bh2587_w60_0_c25 :  std_logic;
signal bh2587_w61_0_c25 :  std_logic;
signal bh2587_w62_0_c25 :  std_logic;
signal bh2587_w63_0_c25 :  std_logic;
signal bh2587_w64_0_c25 :  std_logic;
signal bh2587_w65_0_c25 :  std_logic;
signal bh2587_w66_0_c25 :  std_logic;
signal bh2587_w67_0_c25 :  std_logic;
signal bh2587_w68_0_c25 :  std_logic;
signal bh2587_w69_0_c25 :  std_logic;
signal tile_1_X_c20 :  std_logic_vector(0 downto 0);
signal tile_1_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_1_output_c24 :  std_logic_vector(0 downto 0);
signal tile_1_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_1_c24, bh2587_w39_1_c25 :  std_logic;
signal tile_2_X_c20 :  std_logic_vector(0 downto 0);
signal tile_2_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_2_output_c24 :  std_logic_vector(0 downto 0);
signal tile_2_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_2_c24, bh2587_w39_2_c25 :  std_logic;
signal tile_3_X_c20 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_3_output_c24 :  std_logic_vector(3 downto 0);
signal tile_3_filtered_output_c24 :  unsigned(3-0 downto 0);
signal bh2587_w39_3_c24, bh2587_w39_3_c25 :  std_logic;
signal bh2587_w40_1_c24 :  std_logic;
signal bh2587_w41_1_c24, bh2587_w41_1_c25 :  std_logic;
signal bh2587_w42_1_c24, bh2587_w42_1_c25 :  std_logic;
signal tile_4_X_c20 :  std_logic_vector(0 downto 0);
signal tile_4_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_4_output_c24 :  std_logic_vector(0 downto 0);
signal tile_4_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_4_c24, bh2587_w39_4_c25 :  std_logic;
signal tile_5_X_c20 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_5_output_c24 :  std_logic_vector(1 downto 0);
signal tile_5_filtered_output_c24 :  unsigned(1-0 downto 0);
signal bh2587_w39_5_c24, bh2587_w39_5_c25 :  std_logic;
signal bh2587_w40_2_c24 :  std_logic;
signal tile_6_X_c20 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_6_output_c24 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w40_3_c24 :  std_logic;
signal bh2587_w41_2_c24, bh2587_w41_2_c25 :  std_logic;
signal bh2587_w42_2_c24, bh2587_w42_2_c25 :  std_logic;
signal bh2587_w43_1_c24 :  std_logic;
signal bh2587_w44_1_c24, bh2587_w44_1_c25 :  std_logic;
signal tile_7_X_c20 :  std_logic_vector(0 downto 0);
signal tile_7_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_7_output_c24 :  std_logic_vector(0 downto 0);
signal tile_7_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_6_c24 :  std_logic;
signal tile_8_X_c20 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_8_output_c24 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w39_7_c24 :  std_logic;
signal bh2587_w40_4_c24 :  std_logic;
signal bh2587_w41_3_c24, bh2587_w41_3_c25 :  std_logic;
signal bh2587_w42_3_c24, bh2587_w42_3_c25 :  std_logic;
signal bh2587_w43_2_c24 :  std_logic;
signal tile_9_X_c20 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_9_output_c24 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w42_4_c24, bh2587_w42_4_c25 :  std_logic;
signal bh2587_w43_3_c24 :  std_logic;
signal bh2587_w44_2_c24, bh2587_w44_2_c25 :  std_logic;
signal bh2587_w45_1_c24, bh2587_w45_1_c25 :  std_logic;
signal bh2587_w46_1_c24, bh2587_w46_1_c25 :  std_logic;
signal tile_10_X_c20 :  std_logic_vector(0 downto 0);
signal tile_10_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_10_output_c24 :  std_logic_vector(0 downto 0);
signal tile_10_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_8_c24 :  std_logic;
signal tile_11_X_c20 :  std_logic_vector(1 downto 0);
signal tile_11_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_11_output_c24 :  std_logic_vector(3 downto 0);
signal tile_11_filtered_output_c24 :  unsigned(3-0 downto 0);
signal bh2587_w39_9_c24 :  std_logic;
signal bh2587_w40_5_c24 :  std_logic;
signal bh2587_w41_4_c24, bh2587_w41_4_c25 :  std_logic;
signal bh2587_w42_5_c24, bh2587_w42_5_c25 :  std_logic;
signal tile_12_X_c20 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_12_output_c24 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w41_5_c24, bh2587_w41_5_c25 :  std_logic;
signal bh2587_w42_6_c24, bh2587_w42_6_c25 :  std_logic;
signal bh2587_w43_4_c24 :  std_logic;
signal bh2587_w44_3_c24, bh2587_w44_3_c25 :  std_logic;
signal bh2587_w45_2_c24, bh2587_w45_2_c25 :  std_logic;
signal tile_13_X_c20 :  std_logic_vector(2 downto 0);
signal tile_13_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_13_output_c24 :  std_logic_vector(4 downto 0);
signal tile_13_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w44_4_c24, bh2587_w44_4_c25 :  std_logic;
signal bh2587_w45_3_c24, bh2587_w45_3_c25 :  std_logic;
signal bh2587_w46_2_c24, bh2587_w46_2_c25 :  std_logic;
signal bh2587_w47_1_c24, bh2587_w47_1_c25 :  std_logic;
signal bh2587_w48_1_c24, bh2587_w48_1_c25 :  std_logic;
signal tile_14_X_c20 :  std_logic_vector(0 downto 0);
signal tile_14_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_14_output_c24 :  std_logic_vector(0 downto 0);
signal tile_14_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_10_c24 :  std_logic;
signal tile_15_X_c20 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_15_output_c24 :  std_logic_vector(1 downto 0);
signal tile_15_filtered_output_c24 :  unsigned(1-0 downto 0);
signal bh2587_w39_11_c24 :  std_logic;
signal bh2587_w40_6_c24, bh2587_w40_6_c25 :  std_logic;
signal tile_16_X_c20 :  std_logic_vector(2 downto 0);
signal tile_16_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_16_output_c24 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w40_7_c24, bh2587_w40_7_c25 :  std_logic;
signal bh2587_w41_6_c24, bh2587_w41_6_c25 :  std_logic;
signal bh2587_w42_7_c24, bh2587_w42_7_c25 :  std_logic;
signal bh2587_w43_5_c24 :  std_logic;
signal bh2587_w44_5_c24, bh2587_w44_5_c25 :  std_logic;
signal tile_17_X_c20 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_17_output_c24 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w43_6_c24, bh2587_w43_6_c25 :  std_logic;
signal bh2587_w44_6_c24, bh2587_w44_6_c25 :  std_logic;
signal bh2587_w45_4_c24, bh2587_w45_4_c25 :  std_logic;
signal bh2587_w46_3_c24, bh2587_w46_3_c25 :  std_logic;
signal bh2587_w47_2_c24, bh2587_w47_2_c25 :  std_logic;
signal tile_18_X_c20 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_18_output_c24 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w46_4_c24, bh2587_w46_4_c25 :  std_logic;
signal bh2587_w47_3_c24, bh2587_w47_3_c25 :  std_logic;
signal bh2587_w48_2_c24, bh2587_w48_2_c25 :  std_logic;
signal bh2587_w49_1_c24, bh2587_w49_1_c25 :  std_logic;
signal bh2587_w50_1_c24, bh2587_w50_1_c25 :  std_logic;
signal tile_19_X_c20 :  std_logic_vector(0 downto 0);
signal tile_19_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_19_output_c24 :  std_logic_vector(0 downto 0);
signal tile_19_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_12_c24 :  std_logic;
signal tile_20_X_c20 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_20_output_c24 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w39_13_c24 :  std_logic;
signal bh2587_w40_8_c24, bh2587_w40_8_c25 :  std_logic;
signal bh2587_w41_7_c24, bh2587_w41_7_c25 :  std_logic;
signal bh2587_w42_8_c24, bh2587_w42_8_c25 :  std_logic;
signal bh2587_w43_7_c24, bh2587_w43_7_c25 :  std_logic;
signal tile_21_X_c20 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_21_output_c24 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w42_9_c24, bh2587_w42_9_c25 :  std_logic;
signal bh2587_w43_8_c24, bh2587_w43_8_c25 :  std_logic;
signal bh2587_w44_7_c24, bh2587_w44_7_c25 :  std_logic;
signal bh2587_w45_5_c24, bh2587_w45_5_c25 :  std_logic;
signal bh2587_w46_5_c24, bh2587_w46_5_c25 :  std_logic;
signal tile_22_X_c20 :  std_logic_vector(2 downto 0);
signal tile_22_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_22_output_c24 :  std_logic_vector(4 downto 0);
signal tile_22_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w45_6_c24, bh2587_w45_6_c25 :  std_logic;
signal bh2587_w46_6_c24, bh2587_w46_6_c25 :  std_logic;
signal bh2587_w47_4_c24, bh2587_w47_4_c25 :  std_logic;
signal bh2587_w48_3_c24, bh2587_w48_3_c25 :  std_logic;
signal bh2587_w49_2_c24, bh2587_w49_2_c25 :  std_logic;
signal tile_23_X_c20 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_23_output_c24 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w48_4_c24, bh2587_w48_4_c25 :  std_logic;
signal bh2587_w49_3_c24, bh2587_w49_3_c25 :  std_logic;
signal bh2587_w50_2_c24, bh2587_w50_2_c25 :  std_logic;
signal bh2587_w51_1_c24, bh2587_w51_1_c25 :  std_logic;
signal bh2587_w52_1_c24, bh2587_w52_1_c25 :  std_logic;
signal tile_24_X_c20 :  std_logic_vector(16 downto 0);
signal tile_24_Y_c24 :  std_logic_vector(22 downto 0);
signal tile_24_output_c25 :  std_logic_vector(39 downto 0);
signal tile_24_filtered_output_c25 :  unsigned(39-0 downto 0);
signal bh2587_w53_1_c25 :  std_logic;
signal bh2587_w54_1_c25 :  std_logic;
signal bh2587_w55_1_c25 :  std_logic;
signal bh2587_w56_1_c25 :  std_logic;
signal bh2587_w57_1_c25 :  std_logic;
signal bh2587_w58_1_c25 :  std_logic;
signal bh2587_w59_1_c25 :  std_logic;
signal bh2587_w60_1_c25 :  std_logic;
signal bh2587_w61_1_c25 :  std_logic;
signal bh2587_w62_1_c25 :  std_logic;
signal bh2587_w63_1_c25 :  std_logic;
signal bh2587_w64_1_c25 :  std_logic;
signal bh2587_w65_1_c25 :  std_logic;
signal bh2587_w66_1_c25 :  std_logic;
signal bh2587_w67_1_c25 :  std_logic;
signal bh2587_w68_1_c25 :  std_logic;
signal bh2587_w69_1_c25 :  std_logic;
signal bh2587_w70_0_c25 :  std_logic;
signal bh2587_w71_0_c25 :  std_logic;
signal bh2587_w72_0_c25 :  std_logic;
signal bh2587_w73_0_c25 :  std_logic;
signal bh2587_w74_0_c25 :  std_logic;
signal bh2587_w75_0_c25 :  std_logic;
signal bh2587_w76_0_c25 :  std_logic;
signal bh2587_w77_0_c25 :  std_logic;
signal bh2587_w78_0_c25 :  std_logic;
signal bh2587_w79_0_c25 :  std_logic;
signal bh2587_w80_0_c25 :  std_logic;
signal bh2587_w81_0_c25 :  std_logic;
signal bh2587_w82_0_c25 :  std_logic;
signal bh2587_w83_0_c25 :  std_logic;
signal bh2587_w84_0_c25, bh2587_w84_0_c26 :  std_logic;
signal bh2587_w85_0_c25, bh2587_w85_0_c26 :  std_logic;
signal bh2587_w86_0_c25, bh2587_w86_0_c26 :  std_logic;
signal bh2587_w87_0_c25, bh2587_w87_0_c26 :  std_logic;
signal bh2587_w88_0_c25, bh2587_w88_0_c26 :  std_logic;
signal bh2587_w89_0_c25, bh2587_w89_0_c26 :  std_logic;
signal bh2587_w90_0_c25, bh2587_w90_0_c26 :  std_logic;
signal bh2587_w91_0_c25, bh2587_w91_0_c26 :  std_logic;
signal bh2587_w92_0_c25, bh2587_w92_0_c26 :  std_logic;
signal tile_25_X_c20 :  std_logic_vector(16 downto 0);
signal tile_25_Y_c24 :  std_logic_vector(22 downto 0);
signal tile_25_output_c25 :  std_logic_vector(39 downto 0);
signal tile_25_filtered_output_c25 :  unsigned(39-0 downto 0);
signal bh2587_w36_1_c25 :  std_logic;
signal bh2587_w37_1_c25 :  std_logic;
signal bh2587_w38_1_c25 :  std_logic;
signal bh2587_w39_14_c25 :  std_logic;
signal bh2587_w40_9_c25 :  std_logic;
signal bh2587_w41_8_c25 :  std_logic;
signal bh2587_w42_10_c25 :  std_logic;
signal bh2587_w43_9_c25 :  std_logic;
signal bh2587_w44_8_c25 :  std_logic;
signal bh2587_w45_7_c25 :  std_logic;
signal bh2587_w46_7_c25 :  std_logic;
signal bh2587_w47_5_c25 :  std_logic;
signal bh2587_w48_5_c25 :  std_logic;
signal bh2587_w49_4_c25 :  std_logic;
signal bh2587_w50_3_c25 :  std_logic;
signal bh2587_w51_2_c25 :  std_logic;
signal bh2587_w52_2_c25 :  std_logic;
signal bh2587_w53_2_c25 :  std_logic;
signal bh2587_w54_2_c25 :  std_logic;
signal bh2587_w55_2_c25 :  std_logic;
signal bh2587_w56_2_c25 :  std_logic;
signal bh2587_w57_2_c25 :  std_logic;
signal bh2587_w58_2_c25 :  std_logic;
signal bh2587_w59_2_c25 :  std_logic;
signal bh2587_w60_2_c25 :  std_logic;
signal bh2587_w61_2_c25 :  std_logic;
signal bh2587_w62_2_c25 :  std_logic;
signal bh2587_w63_2_c25 :  std_logic;
signal bh2587_w64_2_c25 :  std_logic;
signal bh2587_w65_2_c25 :  std_logic;
signal bh2587_w66_2_c25 :  std_logic;
signal bh2587_w67_2_c25 :  std_logic;
signal bh2587_w68_2_c25 :  std_logic;
signal bh2587_w69_2_c25 :  std_logic;
signal bh2587_w70_1_c25 :  std_logic;
signal bh2587_w71_1_c25 :  std_logic;
signal bh2587_w72_1_c25 :  std_logic;
signal bh2587_w73_1_c25 :  std_logic;
signal bh2587_w74_1_c25 :  std_logic;
signal bh2587_w75_1_c25 :  std_logic;
signal tile_26_X_c20 :  std_logic_vector(0 downto 0);
signal tile_26_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_26_output_c24 :  std_logic_vector(0 downto 0);
signal tile_26_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_15_c24 :  std_logic;
signal tile_27_X_c20 :  std_logic_vector(0 downto 0);
signal tile_27_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_27_output_c24 :  std_logic_vector(0 downto 0);
signal tile_27_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_16_c24 :  std_logic;
signal tile_28_X_c20 :  std_logic_vector(1 downto 0);
signal tile_28_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_28_output_c24 :  std_logic_vector(3 downto 0);
signal tile_28_filtered_output_c24 :  unsigned(3-0 downto 0);
signal bh2587_w39_17_c24 :  std_logic;
signal bh2587_w40_10_c24 :  std_logic;
signal bh2587_w41_9_c24 :  std_logic;
signal bh2587_w42_11_c24 :  std_logic;
signal tile_29_X_c20 :  std_logic_vector(0 downto 0);
signal tile_29_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_29_output_c24 :  std_logic_vector(0 downto 0);
signal tile_29_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_18_c24 :  std_logic;
signal tile_30_X_c20 :  std_logic_vector(1 downto 0);
signal tile_30_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_30_output_c24 :  std_logic_vector(1 downto 0);
signal tile_30_filtered_output_c24 :  unsigned(1-0 downto 0);
signal bh2587_w39_19_c24 :  std_logic;
signal bh2587_w40_11_c24, bh2587_w40_11_c25 :  std_logic;
signal tile_31_X_c20 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_31_output_c24 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w40_12_c24, bh2587_w40_12_c25 :  std_logic;
signal bh2587_w41_10_c24, bh2587_w41_10_c25 :  std_logic;
signal bh2587_w42_12_c24, bh2587_w42_12_c25 :  std_logic;
signal bh2587_w43_10_c24 :  std_logic;
signal bh2587_w44_9_c24, bh2587_w44_9_c25 :  std_logic;
signal tile_32_X_c20 :  std_logic_vector(0 downto 0);
signal tile_32_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_32_output_c24 :  std_logic_vector(0 downto 0);
signal tile_32_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_20_c24 :  std_logic;
signal tile_33_X_c20 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_33_output_c24 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w39_21_c24 :  std_logic;
signal bh2587_w40_13_c24 :  std_logic;
signal bh2587_w41_11_c24, bh2587_w41_11_c25 :  std_logic;
signal bh2587_w42_13_c24 :  std_logic;
signal bh2587_w43_11_c24 :  std_logic;
signal tile_34_X_c20 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_34_output_c24 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w42_14_c24 :  std_logic;
signal bh2587_w43_12_c24, bh2587_w43_12_c25 :  std_logic;
signal bh2587_w44_10_c24 :  std_logic;
signal bh2587_w45_8_c24, bh2587_w45_8_c25 :  std_logic;
signal bh2587_w46_8_c24, bh2587_w46_8_c25 :  std_logic;
signal tile_35_X_c20 :  std_logic_vector(0 downto 0);
signal tile_35_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_35_output_c24 :  std_logic_vector(0 downto 0);
signal tile_35_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_22_c24 :  std_logic;
signal tile_36_X_c20 :  std_logic_vector(1 downto 0);
signal tile_36_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_36_output_c24 :  std_logic_vector(3 downto 0);
signal tile_36_filtered_output_c24 :  unsigned(3-0 downto 0);
signal bh2587_w39_23_c24, bh2587_w39_23_c25 :  std_logic;
signal bh2587_w40_14_c24 :  std_logic;
signal bh2587_w41_12_c24, bh2587_w41_12_c25 :  std_logic;
signal bh2587_w42_15_c24 :  std_logic;
signal tile_37_X_c20 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_37_output_c24 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w41_13_c24 :  std_logic;
signal bh2587_w42_16_c24 :  std_logic;
signal bh2587_w43_13_c24 :  std_logic;
signal bh2587_w44_11_c24, bh2587_w44_11_c25 :  std_logic;
signal bh2587_w45_9_c24 :  std_logic;
signal tile_38_X_c20 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_38_output_c24 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w44_12_c24, bh2587_w44_12_c25 :  std_logic;
signal bh2587_w45_10_c24, bh2587_w45_10_c25 :  std_logic;
signal bh2587_w46_9_c24 :  std_logic;
signal bh2587_w47_6_c24 :  std_logic;
signal bh2587_w48_6_c24, bh2587_w48_6_c25 :  std_logic;
signal tile_39_X_c20 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_39_output_c24 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c24 :  unsigned(0-0 downto 0);
signal bh2587_w39_24_c24, bh2587_w39_24_c25 :  std_logic;
signal tile_40_X_c20 :  std_logic_vector(1 downto 0);
signal tile_40_Y_c24 :  std_logic_vector(0 downto 0);
signal tile_40_output_c24 :  std_logic_vector(1 downto 0);
signal tile_40_filtered_output_c24 :  unsigned(1-0 downto 0);
signal bh2587_w39_25_c24, bh2587_w39_25_c25 :  std_logic;
signal bh2587_w40_15_c24 :  std_logic;
signal tile_41_X_c20 :  std_logic_vector(2 downto 0);
signal tile_41_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_41_output_c24 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w40_16_c24 :  std_logic;
signal bh2587_w41_14_c24 :  std_logic;
signal bh2587_w42_17_c24 :  std_logic;
signal bh2587_w43_14_c24 :  std_logic;
signal bh2587_w44_13_c24 :  std_logic;
signal tile_42_X_c20 :  std_logic_vector(2 downto 0);
signal tile_42_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_42_output_c24 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w43_15_c24 :  std_logic;
signal bh2587_w44_14_c24 :  std_logic;
signal bh2587_w45_11_c24, bh2587_w45_11_c25 :  std_logic;
signal bh2587_w46_10_c24, bh2587_w46_10_c25 :  std_logic;
signal bh2587_w47_7_c24 :  std_logic;
signal tile_43_X_c20 :  std_logic_vector(2 downto 0);
signal tile_43_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_43_output_c24 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w46_11_c24, bh2587_w46_11_c25 :  std_logic;
signal bh2587_w47_8_c24 :  std_logic;
signal bh2587_w48_7_c24, bh2587_w48_7_c25 :  std_logic;
signal bh2587_w49_5_c24, bh2587_w49_5_c25 :  std_logic;
signal bh2587_w50_4_c24 :  std_logic;
signal tile_44_X_c20 :  std_logic_vector(2 downto 0);
signal tile_44_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_44_output_c24 :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w39_26_c24, bh2587_w39_26_c25 :  std_logic;
signal bh2587_w40_17_c24 :  std_logic;
signal bh2587_w41_15_c24 :  std_logic;
signal bh2587_w42_18_c24 :  std_logic;
signal bh2587_w43_16_c24 :  std_logic;
signal tile_45_X_c20 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_45_output_c24 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w42_19_c24 :  std_logic;
signal bh2587_w43_17_c24 :  std_logic;
signal bh2587_w44_15_c24 :  std_logic;
signal bh2587_w45_12_c24, bh2587_w45_12_c25 :  std_logic;
signal bh2587_w46_12_c24, bh2587_w46_12_c25 :  std_logic;
signal tile_46_X_c20 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_46_output_c24 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w45_13_c24 :  std_logic;
signal bh2587_w46_13_c24 :  std_logic;
signal bh2587_w47_9_c24 :  std_logic;
signal bh2587_w48_8_c24 :  std_logic;
signal bh2587_w49_6_c24, bh2587_w49_6_c25 :  std_logic;
signal tile_47_X_c20 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_47_output_c24 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w48_9_c24, bh2587_w48_9_c25 :  std_logic;
signal bh2587_w49_7_c24 :  std_logic;
signal bh2587_w50_5_c24 :  std_logic;
signal bh2587_w51_3_c24 :  std_logic;
signal bh2587_w52_3_c24, bh2587_w52_3_c25 :  std_logic;
signal tile_48_X_c20 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_48_output_c24 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w41_16_c24 :  std_logic;
signal bh2587_w42_20_c24 :  std_logic;
signal bh2587_w43_18_c24 :  std_logic;
signal bh2587_w44_16_c24 :  std_logic;
signal bh2587_w45_14_c24 :  std_logic;
signal tile_49_X_c20 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_49_output_c24 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w44_17_c24 :  std_logic;
signal bh2587_w45_15_c24 :  std_logic;
signal bh2587_w46_14_c24 :  std_logic;
signal bh2587_w47_10_c24 :  std_logic;
signal bh2587_w48_10_c24 :  std_logic;
signal tile_50_X_c20 :  std_logic_vector(2 downto 0);
signal tile_50_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_50_output_c24 :  std_logic_vector(4 downto 0);
signal tile_50_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w47_11_c24 :  std_logic;
signal bh2587_w48_11_c24 :  std_logic;
signal bh2587_w49_8_c24 :  std_logic;
signal bh2587_w50_6_c24 :  std_logic;
signal bh2587_w51_4_c24 :  std_logic;
signal tile_51_X_c20 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_51_output_c24 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w50_7_c24 :  std_logic;
signal bh2587_w51_5_c24 :  std_logic;
signal bh2587_w52_4_c24, bh2587_w52_4_c25 :  std_logic;
signal bh2587_w53_3_c24, bh2587_w53_3_c25 :  std_logic;
signal bh2587_w54_3_c24, bh2587_w54_3_c25 :  std_logic;
signal tile_52_X_c20 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_52_output_c24 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w43_19_c24 :  std_logic;
signal bh2587_w44_18_c24 :  std_logic;
signal bh2587_w45_16_c24 :  std_logic;
signal bh2587_w46_15_c24 :  std_logic;
signal bh2587_w47_12_c24 :  std_logic;
signal tile_53_X_c20 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_53_output_c24 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w46_16_c24 :  std_logic;
signal bh2587_w47_13_c24 :  std_logic;
signal bh2587_w48_12_c24 :  std_logic;
signal bh2587_w49_9_c24 :  std_logic;
signal bh2587_w50_8_c24 :  std_logic;
signal tile_54_X_c20 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_54_output_c24 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w49_10_c24 :  std_logic;
signal bh2587_w50_9_c24 :  std_logic;
signal bh2587_w51_6_c24 :  std_logic;
signal bh2587_w52_5_c24, bh2587_w52_5_c25 :  std_logic;
signal bh2587_w53_4_c24, bh2587_w53_4_c25 :  std_logic;
signal tile_55_X_c20 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_55_output_c24 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w52_6_c24 :  std_logic;
signal bh2587_w53_5_c24, bh2587_w53_5_c25 :  std_logic;
signal bh2587_w54_4_c24, bh2587_w54_4_c25 :  std_logic;
signal bh2587_w55_3_c24, bh2587_w55_3_c25 :  std_logic;
signal bh2587_w56_3_c24, bh2587_w56_3_c25 :  std_logic;
signal tile_56_X_c20 :  std_logic_vector(2 downto 0);
signal tile_56_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_56_output_c24 :  std_logic_vector(4 downto 0);
signal tile_56_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w45_17_c24 :  std_logic;
signal bh2587_w46_17_c24 :  std_logic;
signal bh2587_w47_14_c24 :  std_logic;
signal bh2587_w48_13_c24 :  std_logic;
signal bh2587_w49_11_c24 :  std_logic;
signal tile_57_X_c20 :  std_logic_vector(2 downto 0);
signal tile_57_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_57_output_c24 :  std_logic_vector(4 downto 0);
signal tile_57_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w48_14_c24 :  std_logic;
signal bh2587_w49_12_c24 :  std_logic;
signal bh2587_w50_10_c24 :  std_logic;
signal bh2587_w51_7_c24 :  std_logic;
signal bh2587_w52_7_c24 :  std_logic;
signal tile_58_X_c20 :  std_logic_vector(2 downto 0);
signal tile_58_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_58_output_c24 :  std_logic_vector(4 downto 0);
signal tile_58_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w51_8_c24 :  std_logic;
signal bh2587_w52_8_c24 :  std_logic;
signal bh2587_w53_6_c24, bh2587_w53_6_c25 :  std_logic;
signal bh2587_w54_5_c24, bh2587_w54_5_c25 :  std_logic;
signal bh2587_w55_4_c24, bh2587_w55_4_c25 :  std_logic;
signal tile_59_X_c20 :  std_logic_vector(2 downto 0);
signal tile_59_Y_c24 :  std_logic_vector(1 downto 0);
signal tile_59_output_c24 :  std_logic_vector(4 downto 0);
signal tile_59_filtered_output_c24 :  unsigned(4-0 downto 0);
signal bh2587_w54_6_c24 :  std_logic;
signal bh2587_w55_5_c24, bh2587_w55_5_c25 :  std_logic;
signal bh2587_w56_4_c24, bh2587_w56_4_c25 :  std_logic;
signal bh2587_w57_3_c24, bh2587_w57_3_c25 :  std_logic;
signal bh2587_w58_3_c24, bh2587_w58_3_c25 :  std_logic;
signal bh2587_w39_27_c0, bh2587_w39_27_c1, bh2587_w39_27_c2, bh2587_w39_27_c3, bh2587_w39_27_c4, bh2587_w39_27_c5, bh2587_w39_27_c6, bh2587_w39_27_c7, bh2587_w39_27_c8, bh2587_w39_27_c9, bh2587_w39_27_c10, bh2587_w39_27_c11, bh2587_w39_27_c12, bh2587_w39_27_c13, bh2587_w39_27_c14, bh2587_w39_27_c15, bh2587_w39_27_c16, bh2587_w39_27_c17, bh2587_w39_27_c18, bh2587_w39_27_c19, bh2587_w39_27_c20, bh2587_w39_27_c21, bh2587_w39_27_c22, bh2587_w39_27_c23, bh2587_w39_27_c24, bh2587_w39_27_c25 :  std_logic;
signal bh2587_w40_18_c0, bh2587_w40_18_c1, bh2587_w40_18_c2, bh2587_w40_18_c3, bh2587_w40_18_c4, bh2587_w40_18_c5, bh2587_w40_18_c6, bh2587_w40_18_c7, bh2587_w40_18_c8, bh2587_w40_18_c9, bh2587_w40_18_c10, bh2587_w40_18_c11, bh2587_w40_18_c12, bh2587_w40_18_c13, bh2587_w40_18_c14, bh2587_w40_18_c15, bh2587_w40_18_c16, bh2587_w40_18_c17, bh2587_w40_18_c18, bh2587_w40_18_c19, bh2587_w40_18_c20, bh2587_w40_18_c21, bh2587_w40_18_c22, bh2587_w40_18_c23, bh2587_w40_18_c24 :  std_logic;
signal bh2587_w41_17_c0, bh2587_w41_17_c1, bh2587_w41_17_c2, bh2587_w41_17_c3, bh2587_w41_17_c4, bh2587_w41_17_c5, bh2587_w41_17_c6, bh2587_w41_17_c7, bh2587_w41_17_c8, bh2587_w41_17_c9, bh2587_w41_17_c10, bh2587_w41_17_c11, bh2587_w41_17_c12, bh2587_w41_17_c13, bh2587_w41_17_c14, bh2587_w41_17_c15, bh2587_w41_17_c16, bh2587_w41_17_c17, bh2587_w41_17_c18, bh2587_w41_17_c19, bh2587_w41_17_c20, bh2587_w41_17_c21, bh2587_w41_17_c22, bh2587_w41_17_c23, bh2587_w41_17_c24 :  std_logic;
signal bh2587_w42_21_c0, bh2587_w42_21_c1, bh2587_w42_21_c2, bh2587_w42_21_c3, bh2587_w42_21_c4, bh2587_w42_21_c5, bh2587_w42_21_c6, bh2587_w42_21_c7, bh2587_w42_21_c8, bh2587_w42_21_c9, bh2587_w42_21_c10, bh2587_w42_21_c11, bh2587_w42_21_c12, bh2587_w42_21_c13, bh2587_w42_21_c14, bh2587_w42_21_c15, bh2587_w42_21_c16, bh2587_w42_21_c17, bh2587_w42_21_c18, bh2587_w42_21_c19, bh2587_w42_21_c20, bh2587_w42_21_c21, bh2587_w42_21_c22, bh2587_w42_21_c23, bh2587_w42_21_c24 :  std_logic;
signal bh2587_w43_20_c0, bh2587_w43_20_c1, bh2587_w43_20_c2, bh2587_w43_20_c3, bh2587_w43_20_c4, bh2587_w43_20_c5, bh2587_w43_20_c6, bh2587_w43_20_c7, bh2587_w43_20_c8, bh2587_w43_20_c9, bh2587_w43_20_c10, bh2587_w43_20_c11, bh2587_w43_20_c12, bh2587_w43_20_c13, bh2587_w43_20_c14, bh2587_w43_20_c15, bh2587_w43_20_c16, bh2587_w43_20_c17, bh2587_w43_20_c18, bh2587_w43_20_c19, bh2587_w43_20_c20, bh2587_w43_20_c21, bh2587_w43_20_c22, bh2587_w43_20_c23, bh2587_w43_20_c24 :  std_logic;
signal bh2587_w44_19_c0, bh2587_w44_19_c1, bh2587_w44_19_c2, bh2587_w44_19_c3, bh2587_w44_19_c4, bh2587_w44_19_c5, bh2587_w44_19_c6, bh2587_w44_19_c7, bh2587_w44_19_c8, bh2587_w44_19_c9, bh2587_w44_19_c10, bh2587_w44_19_c11, bh2587_w44_19_c12, bh2587_w44_19_c13, bh2587_w44_19_c14, bh2587_w44_19_c15, bh2587_w44_19_c16, bh2587_w44_19_c17, bh2587_w44_19_c18, bh2587_w44_19_c19, bh2587_w44_19_c20, bh2587_w44_19_c21, bh2587_w44_19_c22, bh2587_w44_19_c23, bh2587_w44_19_c24 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2831_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2831_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w36_2_c25, bh2587_w36_2_c26 :  std_logic;
signal bh2587_w37_2_c25 :  std_logic;
signal bh2587_w38_2_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_copy2832_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2835_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w38_3_c25 :  std_logic;
signal bh2587_w39_28_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_copy2836_c25 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2839_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w39_29_c25 :  std_logic;
signal bh2587_w40_19_c25 :  std_logic;
signal bh2587_w41_18_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_copy2840_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2841_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w39_30_c25 :  std_logic;
signal bh2587_w40_20_c25 :  std_logic;
signal bh2587_w41_19_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_copy2842_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2843_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w39_31_c24, bh2587_w39_31_c25 :  std_logic;
signal bh2587_w40_21_c24, bh2587_w40_21_c25 :  std_logic;
signal bh2587_w41_20_c24, bh2587_w41_20_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_copy2844_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2845_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w39_32_c24, bh2587_w39_32_c25 :  std_logic;
signal bh2587_w40_22_c24, bh2587_w40_22_c25 :  std_logic;
signal bh2587_w41_21_c24, bh2587_w41_21_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_copy2846_c24 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In0_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w39_33_c25 :  std_logic;
signal bh2587_w40_23_c25 :  std_logic;
signal bh2587_w41_22_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_copy2850_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2851_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w40_24_c24, bh2587_w40_24_c25 :  std_logic;
signal bh2587_w41_23_c24, bh2587_w41_23_c25 :  std_logic;
signal bh2587_w42_22_c24, bh2587_w42_22_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_copy2852_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2853_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w40_25_c24, bh2587_w40_25_c25 :  std_logic;
signal bh2587_w41_24_c24, bh2587_w41_24_c25 :  std_logic;
signal bh2587_w42_23_c24, bh2587_w42_23_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_copy2854_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2855_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w40_26_c25 :  std_logic;
signal bh2587_w41_25_c25 :  std_logic;
signal bh2587_w42_24_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_copy2856_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2857_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w41_26_c24, bh2587_w41_26_c25 :  std_logic;
signal bh2587_w42_25_c24, bh2587_w42_25_c25 :  std_logic;
signal bh2587_w43_21_c24, bh2587_w43_21_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_copy2858_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2859_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w41_27_c25 :  std_logic;
signal bh2587_w42_26_c25 :  std_logic;
signal bh2587_w43_22_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_copy2860_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2861_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w41_28_c25 :  std_logic;
signal bh2587_w42_27_c25 :  std_logic;
signal bh2587_w43_23_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_copy2862_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2863_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w42_28_c25 :  std_logic;
signal bh2587_w43_24_c25 :  std_logic;
signal bh2587_w44_20_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_copy2864_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2865_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w42_29_c24, bh2587_w42_29_c25 :  std_logic;
signal bh2587_w43_25_c24, bh2587_w43_25_c25 :  std_logic;
signal bh2587_w44_21_c24, bh2587_w44_21_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_copy2866_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2867_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w42_30_c25 :  std_logic;
signal bh2587_w43_26_c25 :  std_logic;
signal bh2587_w44_22_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_copy2868_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In0_c24 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c24 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w42_31_c24, bh2587_w42_31_c25 :  std_logic;
signal bh2587_w43_27_c24, bh2587_w43_27_c25 :  std_logic;
signal bh2587_w44_23_c24 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_copy2870_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2871_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w43_28_c24, bh2587_w43_28_c25 :  std_logic;
signal bh2587_w44_24_c24, bh2587_w44_24_c25 :  std_logic;
signal bh2587_w45_18_c24, bh2587_w45_18_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_copy2872_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2873_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w43_29_c24, bh2587_w43_29_c25 :  std_logic;
signal bh2587_w44_25_c24 :  std_logic;
signal bh2587_w45_19_c24, bh2587_w45_19_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_copy2874_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2875_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w43_30_c25 :  std_logic;
signal bh2587_w44_26_c25 :  std_logic;
signal bh2587_w45_20_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_copy2876_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2877_In0_c24 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2877_In1_c24 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w43_31_c24, bh2587_w43_31_c25 :  std_logic;
signal bh2587_w44_27_c24 :  std_logic;
signal bh2587_w45_21_c24, bh2587_w45_21_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_copy2878_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2879_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w44_28_c25 :  std_logic;
signal bh2587_w45_22_c25 :  std_logic;
signal bh2587_w46_18_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_copy2880_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2881_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w44_29_c24 :  std_logic;
signal bh2587_w45_23_c24, bh2587_w45_23_c25 :  std_logic;
signal bh2587_w46_19_c24, bh2587_w46_19_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_copy2882_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2883_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w44_30_c25 :  std_logic;
signal bh2587_w45_24_c25 :  std_logic;
signal bh2587_w46_20_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_copy2884_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2885_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w45_25_c24, bh2587_w45_25_c25 :  std_logic;
signal bh2587_w46_21_c24, bh2587_w46_21_c25 :  std_logic;
signal bh2587_w47_15_c24, bh2587_w47_15_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_copy2886_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2887_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w45_26_c25 :  std_logic;
signal bh2587_w46_22_c25 :  std_logic;
signal bh2587_w47_16_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_copy2888_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2889_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w45_27_c25 :  std_logic;
signal bh2587_w46_23_c25 :  std_logic;
signal bh2587_w47_17_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_copy2890_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2891_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w46_24_c25 :  std_logic;
signal bh2587_w47_18_c25 :  std_logic;
signal bh2587_w48_15_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_copy2892_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2893_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w46_25_c24, bh2587_w46_25_c25 :  std_logic;
signal bh2587_w47_19_c24, bh2587_w47_19_c25 :  std_logic;
signal bh2587_w48_16_c24, bh2587_w48_16_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_copy2894_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2895_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w46_26_c25 :  std_logic;
signal bh2587_w47_20_c25 :  std_logic;
signal bh2587_w48_17_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_copy2896_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2897_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w47_21_c24, bh2587_w47_21_c25 :  std_logic;
signal bh2587_w48_18_c24, bh2587_w48_18_c25 :  std_logic;
signal bh2587_w49_13_c24, bh2587_w49_13_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_copy2898_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2899_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w47_22_c25 :  std_logic;
signal bh2587_w48_19_c25 :  std_logic;
signal bh2587_w49_14_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_copy2900_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In0_c24, Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w47_23_c25 :  std_logic;
signal bh2587_w48_20_c25 :  std_logic;
signal bh2587_w49_15_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_copy2902_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2903_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w48_21_c24, bh2587_w48_21_c25 :  std_logic;
signal bh2587_w49_16_c24, bh2587_w49_16_c25 :  std_logic;
signal bh2587_w50_11_c24, bh2587_w50_11_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_copy2904_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2905_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w48_22_c25 :  std_logic;
signal bh2587_w49_17_c25 :  std_logic;
signal bh2587_w50_12_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_copy2906_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2907_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w49_18_c25 :  std_logic;
signal bh2587_w50_13_c25 :  std_logic;
signal bh2587_w51_9_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_copy2908_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2909_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w49_19_c24, bh2587_w49_19_c25 :  std_logic;
signal bh2587_w50_14_c24, bh2587_w50_14_c25 :  std_logic;
signal bh2587_w51_10_c24, bh2587_w51_10_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_copy2910_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2911_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w50_15_c25 :  std_logic;
signal bh2587_w51_11_c25 :  std_logic;
signal bh2587_w52_9_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_copy2912_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In0_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w50_16_c25 :  std_logic;
signal bh2587_w51_12_c25 :  std_logic;
signal bh2587_w52_10_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_copy2914_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In0_c24, Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w50_17_c25 :  std_logic;
signal bh2587_w51_13_c25 :  std_logic;
signal bh2587_w52_11_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_copy2916_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2917_In0_c24 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_c24 :  std_logic_vector(2 downto 0);
signal bh2587_w51_14_c24, bh2587_w51_14_c25 :  std_logic;
signal bh2587_w52_12_c24, bh2587_w52_12_c25 :  std_logic;
signal bh2587_w53_7_c24, bh2587_w53_7_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_copy2918_c24 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2919_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w52_13_c25 :  std_logic;
signal bh2587_w53_8_c25 :  std_logic;
signal bh2587_w54_7_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_copy2920_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2921_In0_c24 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_c24 :  std_logic_vector(1 downto 0);
signal bh2587_w52_14_c24, bh2587_w52_14_c25 :  std_logic;
signal bh2587_w53_9_c24, bh2587_w53_9_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_copy2922_c24 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2923_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w53_10_c25 :  std_logic;
signal bh2587_w54_8_c25 :  std_logic;
signal bh2587_w55_6_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_copy2924_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2925_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w54_9_c25 :  std_logic;
signal bh2587_w55_7_c25 :  std_logic;
signal bh2587_w56_5_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_copy2926_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2927_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w55_8_c25 :  std_logic;
signal bh2587_w56_6_c25 :  std_logic;
signal bh2587_w57_4_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_copy2928_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2929_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2929_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w56_7_c25 :  std_logic;
signal bh2587_w57_5_c25 :  std_logic;
signal bh2587_w58_4_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_copy2930_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2931_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w57_6_c25 :  std_logic;
signal bh2587_w58_5_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_copy2932_c25 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w58_6_c25 :  std_logic;
signal bh2587_w59_3_c25 :  std_logic;
signal bh2587_w60_3_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_copy2934_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2935_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w59_4_c25 :  std_logic;
signal bh2587_w60_4_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_copy2936_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2937_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2937_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w60_5_c25 :  std_logic;
signal bh2587_w61_3_c25 :  std_logic;
signal bh2587_w62_3_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_copy2938_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2939_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2939_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w62_4_c25 :  std_logic;
signal bh2587_w63_3_c25 :  std_logic;
signal bh2587_w64_3_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_copy2940_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2941_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2941_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w64_4_c25 :  std_logic;
signal bh2587_w65_3_c25 :  std_logic;
signal bh2587_w66_3_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_copy2942_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2943_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2943_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w66_4_c25 :  std_logic;
signal bh2587_w67_3_c25 :  std_logic;
signal bh2587_w68_3_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_copy2944_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2945_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2945_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w68_4_c25 :  std_logic;
signal bh2587_w69_3_c25 :  std_logic;
signal bh2587_w70_2_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_copy2946_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2947_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2947_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w70_3_c25 :  std_logic;
signal bh2587_w71_2_c25 :  std_logic;
signal bh2587_w72_2_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_copy2948_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2949_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2949_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w72_3_c25 :  std_logic;
signal bh2587_w73_2_c25 :  std_logic;
signal bh2587_w74_2_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_copy2950_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2951_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2951_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w74_3_c25 :  std_logic;
signal bh2587_w75_2_c25 :  std_logic;
signal bh2587_w76_1_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_copy2952_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2953_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2953_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w37_3_c25, bh2587_w37_3_c26 :  std_logic;
signal bh2587_w38_4_c25 :  std_logic;
signal bh2587_w39_34_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_copy2954_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2955_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w39_35_c25 :  std_logic;
signal bh2587_w40_27_c25 :  std_logic;
signal bh2587_w41_29_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_copy2956_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2957_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w40_28_c25 :  std_logic;
signal bh2587_w41_30_c25 :  std_logic;
signal bh2587_w42_32_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_copy2958_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2959_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2959_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w40_29_c25 :  std_logic;
signal bh2587_w41_31_c25 :  std_logic;
signal bh2587_w42_33_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_copy2960_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2961_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w41_32_c25 :  std_logic;
signal bh2587_w42_34_c25 :  std_logic;
signal bh2587_w43_32_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_copy2962_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2963_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2963_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w41_33_c25 :  std_logic;
signal bh2587_w42_35_c25 :  std_logic;
signal bh2587_w43_33_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_copy2964_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2965_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w42_36_c25 :  std_logic;
signal bh2587_w43_34_c25 :  std_logic;
signal bh2587_w44_31_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_copy2966_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2967_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w42_37_c25 :  std_logic;
signal bh2587_w43_35_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_copy2968_c25 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2969_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w43_36_c25 :  std_logic;
signal bh2587_w44_32_c25 :  std_logic;
signal bh2587_w45_28_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_copy2970_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2971_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2971_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w43_37_c25 :  std_logic;
signal bh2587_w44_33_c25 :  std_logic;
signal bh2587_w45_29_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_copy2972_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2973_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w44_34_c25 :  std_logic;
signal bh2587_w45_30_c25 :  std_logic;
signal bh2587_w46_27_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_copy2974_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In0_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w44_35_c25 :  std_logic;
signal bh2587_w45_31_c25 :  std_logic;
signal bh2587_w46_28_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_copy2976_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2977_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w45_32_c25 :  std_logic;
signal bh2587_w46_29_c25 :  std_logic;
signal bh2587_w47_24_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_copy2978_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2979_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2979_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w45_33_c25 :  std_logic;
signal bh2587_w46_30_c25 :  std_logic;
signal bh2587_w47_25_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_copy2980_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2981_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w46_31_c25 :  std_logic;
signal bh2587_w47_26_c25 :  std_logic;
signal bh2587_w48_23_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_copy2982_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2983_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w47_27_c25 :  std_logic;
signal bh2587_w48_24_c25 :  std_logic;
signal bh2587_w49_20_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_copy2984_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2985_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2985_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w47_28_c25 :  std_logic;
signal bh2587_w48_25_c25 :  std_logic;
signal bh2587_w49_21_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_copy2986_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2987_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w48_26_c25 :  std_logic;
signal bh2587_w49_22_c25 :  std_logic;
signal bh2587_w50_18_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_copy2988_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2989_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w49_23_c25 :  std_logic;
signal bh2587_w50_19_c25 :  std_logic;
signal bh2587_w51_15_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_copy2990_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2991_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2991_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w49_24_c25 :  std_logic;
signal bh2587_w50_20_c25 :  std_logic;
signal bh2587_w51_16_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_copy2992_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2993_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w50_21_c25 :  std_logic;
signal bh2587_w51_17_c25 :  std_logic;
signal bh2587_w52_15_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_copy2994_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2995_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w51_18_c25 :  std_logic;
signal bh2587_w52_16_c25 :  std_logic;
signal bh2587_w53_11_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_copy2996_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2997_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w52_17_c25 :  std_logic;
signal bh2587_w53_12_c25 :  std_logic;
signal bh2587_w54_10_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_copy2998_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w53_13_c25 :  std_logic;
signal bh2587_w54_11_c25 :  std_logic;
signal bh2587_w55_9_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_copy3000_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3001_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3001_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w54_12_c25 :  std_logic;
signal bh2587_w55_10_c25 :  std_logic;
signal bh2587_w56_8_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_copy3002_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w56_9_c25 :  std_logic;
signal bh2587_w57_7_c25 :  std_logic;
signal bh2587_w58_7_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_copy3004_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3005_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w57_8_c25 :  std_logic;
signal bh2587_w58_8_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_copy3006_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3007_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3007_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w58_9_c25 :  std_logic;
signal bh2587_w59_5_c25 :  std_logic;
signal bh2587_w60_6_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_copy3008_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3009_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3009_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w60_7_c25 :  std_logic;
signal bh2587_w61_4_c25 :  std_logic;
signal bh2587_w62_5_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_copy3010_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3011_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3011_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w62_6_c25 :  std_logic;
signal bh2587_w63_4_c25 :  std_logic;
signal bh2587_w64_5_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_copy3012_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3013_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3013_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w64_6_c25 :  std_logic;
signal bh2587_w65_4_c25 :  std_logic;
signal bh2587_w66_5_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_copy3014_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3015_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3015_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w66_6_c25 :  std_logic;
signal bh2587_w67_4_c25 :  std_logic;
signal bh2587_w68_5_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_copy3016_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3017_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3017_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w68_6_c25 :  std_logic;
signal bh2587_w69_4_c25 :  std_logic;
signal bh2587_w70_4_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_copy3018_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3019_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3019_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w70_5_c25 :  std_logic;
signal bh2587_w71_3_c25 :  std_logic;
signal bh2587_w72_4_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_copy3020_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3021_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3021_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w72_5_c25 :  std_logic;
signal bh2587_w73_3_c25 :  std_logic;
signal bh2587_w74_4_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_copy3022_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3023_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3023_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w74_5_c25 :  std_logic;
signal bh2587_w75_3_c25 :  std_logic;
signal bh2587_w76_2_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_copy3024_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3025_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3025_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w76_3_c25 :  std_logic;
signal bh2587_w77_1_c25 :  std_logic;
signal bh2587_w78_1_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_copy3026_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3027_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3027_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w38_5_c25, bh2587_w38_5_c26 :  std_logic;
signal bh2587_w39_36_c25, bh2587_w39_36_c26 :  std_logic;
signal bh2587_w40_30_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_copy3028_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3029_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w40_31_c25 :  std_logic;
signal bh2587_w41_34_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_copy3030_c25 :  std_logic_vector(1 downto 0);
signal Compressor_5_3_Freq300_uid3032_bh2587_uid3033_In0_c25 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w41_35_c25 :  std_logic;
signal bh2587_w42_38_c25 :  std_logic;
signal bh2587_w43_38_c25 :  std_logic;
signal Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_copy3034_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3035_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w42_39_c25 :  std_logic;
signal bh2587_w43_39_c25 :  std_logic;
signal bh2587_w44_36_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_copy3036_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3037_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w43_40_c25 :  std_logic;
signal bh2587_w44_37_c25 :  std_logic;
signal bh2587_w45_34_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_copy3038_c25 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid3032_bh2587_uid3039_In0_c25 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w44_38_c25 :  std_logic;
signal bh2587_w45_35_c25 :  std_logic;
signal bh2587_w46_32_c25 :  std_logic;
signal Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_copy3040_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3041_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w45_36_c25 :  std_logic;
signal bh2587_w46_33_c25 :  std_logic;
signal bh2587_w47_29_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_copy3042_c25 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3043_In0_c25 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w46_34_c25 :  std_logic;
signal bh2587_w47_30_c25 :  std_logic;
signal bh2587_w48_27_c25 :  std_logic;
signal Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_copy3044_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3045_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3045_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w47_31_c25 :  std_logic;
signal bh2587_w48_28_c25 :  std_logic;
signal bh2587_w49_25_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_copy3046_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3047_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3047_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w48_29_c25 :  std_logic;
signal bh2587_w49_26_c25 :  std_logic;
signal bh2587_w50_22_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_copy3048_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3049_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3049_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w49_27_c25 :  std_logic;
signal bh2587_w50_23_c25 :  std_logic;
signal bh2587_w51_19_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_copy3050_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3051_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w50_24_c25 :  std_logic;
signal bh2587_w51_20_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_copy3052_c25 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w51_21_c25 :  std_logic;
signal bh2587_w52_18_c25 :  std_logic;
signal bh2587_w53_14_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_copy3054_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3055_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w52_19_c25 :  std_logic;
signal bh2587_w53_15_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_copy3056_c25 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w53_16_c25 :  std_logic;
signal bh2587_w54_13_c25 :  std_logic;
signal bh2587_w55_11_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_copy3058_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3059_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w54_14_c25 :  std_logic;
signal bh2587_w55_12_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_copy3060_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3061_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3061_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w55_13_c25 :  std_logic;
signal bh2587_w56_10_c25 :  std_logic;
signal bh2587_w57_9_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_copy3062_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3063_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w57_10_c25 :  std_logic;
signal bh2587_w58_10_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_copy3064_c25 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3065_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w58_11_c25 :  std_logic;
signal bh2587_w59_6_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_copy3066_c25 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3067_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3067_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w60_8_c25 :  std_logic;
signal bh2587_w61_5_c25 :  std_logic;
signal bh2587_w62_7_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_copy3068_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3069_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3069_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w62_8_c25 :  std_logic;
signal bh2587_w63_5_c25 :  std_logic;
signal bh2587_w64_7_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_copy3070_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3071_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3071_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w64_8_c25 :  std_logic;
signal bh2587_w65_5_c25 :  std_logic;
signal bh2587_w66_7_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_copy3072_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3073_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3073_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w66_8_c25 :  std_logic;
signal bh2587_w67_5_c25 :  std_logic;
signal bh2587_w68_7_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_copy3074_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3075_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3075_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w68_8_c25 :  std_logic;
signal bh2587_w69_5_c25 :  std_logic;
signal bh2587_w70_6_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_copy3076_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3077_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3077_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w70_7_c25 :  std_logic;
signal bh2587_w71_4_c25 :  std_logic;
signal bh2587_w72_6_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_copy3078_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3079_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3079_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w72_7_c25 :  std_logic;
signal bh2587_w73_4_c25 :  std_logic;
signal bh2587_w74_6_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_copy3080_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3081_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3081_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w74_7_c25 :  std_logic;
signal bh2587_w75_4_c25 :  std_logic;
signal bh2587_w76_4_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_copy3082_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3083_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3083_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w76_5_c25 :  std_logic;
signal bh2587_w77_2_c25 :  std_logic;
signal bh2587_w78_2_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_copy3084_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3085_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3085_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w78_3_c25 :  std_logic;
signal bh2587_w79_1_c25 :  std_logic;
signal bh2587_w80_1_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_copy3086_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3087_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3087_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w40_32_c25, bh2587_w40_32_c26 :  std_logic;
signal bh2587_w41_36_c25, bh2587_w41_36_c26 :  std_logic;
signal bh2587_w42_40_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_copy3088_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3089_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w42_41_c25 :  std_logic;
signal bh2587_w43_41_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_copy3090_c25 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w43_42_c25 :  std_logic;
signal bh2587_w44_39_c25 :  std_logic;
signal bh2587_w45_37_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_copy3092_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3093_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w44_40_c25 :  std_logic;
signal bh2587_w45_38_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_copy3094_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3095_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3095_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w45_39_c25 :  std_logic;
signal bh2587_w46_35_c25 :  std_logic;
signal bh2587_w47_32_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_copy3096_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c0, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c1, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c2, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c3, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c4, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c5, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c6, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c7, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c8, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c9, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c10, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c11, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c12, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c13, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c14, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c15, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c16, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c17, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c18, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c19, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c20, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c21, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c22, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c23, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c24, Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w47_33_c25 :  std_logic;
signal bh2587_w48_30_c25 :  std_logic;
signal bh2587_w49_28_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_copy3098_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3099_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w48_31_c25 :  std_logic;
signal bh2587_w49_29_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_copy3100_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3101_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3101_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w49_30_c25 :  std_logic;
signal bh2587_w50_25_c25 :  std_logic;
signal bh2587_w51_22_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_copy3102_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3103_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3103_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w51_23_c25 :  std_logic;
signal bh2587_w52_20_c25 :  std_logic;
signal bh2587_w53_17_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_copy3104_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3105_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3105_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w53_18_c25 :  std_logic;
signal bh2587_w54_15_c25 :  std_logic;
signal bh2587_w55_14_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_copy3106_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3107_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_c25 :  std_logic_vector(1 downto 0);
signal bh2587_w55_15_c25 :  std_logic;
signal bh2587_w56_11_c25 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_copy3108_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3109_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3109_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w57_11_c25, bh2587_w57_11_c26 :  std_logic;
signal bh2587_w58_12_c25, bh2587_w58_12_c26 :  std_logic;
signal bh2587_w59_7_c25 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_copy3110_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3111_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3111_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w59_8_c25 :  std_logic;
signal bh2587_w60_9_c25 :  std_logic;
signal bh2587_w61_6_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_copy3112_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3113_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3113_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w62_9_c25 :  std_logic;
signal bh2587_w63_6_c25, bh2587_w63_6_c26 :  std_logic;
signal bh2587_w64_9_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_copy3114_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3115_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3115_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w64_10_c25 :  std_logic;
signal bh2587_w65_6_c25 :  std_logic;
signal bh2587_w66_9_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_copy3116_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3117_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3117_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w66_10_c25 :  std_logic;
signal bh2587_w67_6_c25 :  std_logic;
signal bh2587_w68_9_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_copy3118_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3119_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3119_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w68_10_c25 :  std_logic;
signal bh2587_w69_6_c25 :  std_logic;
signal bh2587_w70_8_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_copy3120_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3121_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3121_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w70_9_c25 :  std_logic;
signal bh2587_w71_5_c25 :  std_logic;
signal bh2587_w72_8_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_copy3122_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3123_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3123_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w72_9_c25 :  std_logic;
signal bh2587_w73_5_c25 :  std_logic;
signal bh2587_w74_8_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_copy3124_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3125_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3125_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w74_9_c25 :  std_logic;
signal bh2587_w75_5_c25 :  std_logic;
signal bh2587_w76_6_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_copy3126_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3127_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3127_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w76_7_c25 :  std_logic;
signal bh2587_w77_3_c25 :  std_logic;
signal bh2587_w78_4_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_copy3128_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3129_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3129_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w78_5_c25 :  std_logic;
signal bh2587_w79_2_c25 :  std_logic;
signal bh2587_w80_2_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_copy3130_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3131_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3131_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w80_3_c25 :  std_logic;
signal bh2587_w81_1_c25 :  std_logic;
signal bh2587_w82_1_c25 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_copy3132_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3133_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3133_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w42_42_c26 :  std_logic;
signal bh2587_w43_43_c26 :  std_logic;
signal bh2587_w44_41_c26 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_copy3134_c25, Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_copy3134_c26 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3135_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_c26 :  std_logic_vector(1 downto 0);
signal bh2587_w44_42_c26 :  std_logic;
signal bh2587_w45_40_c26 :  std_logic;
signal Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_copy3136_c25, Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_copy3136_c26 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3137_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3137_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w45_41_c26 :  std_logic;
signal bh2587_w46_36_c26 :  std_logic;
signal bh2587_w47_34_c26 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_copy3138_c25, Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_copy3138_c26 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3139_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3139_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w47_35_c26 :  std_logic;
signal bh2587_w48_32_c26 :  std_logic;
signal bh2587_w49_31_c26 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_copy3140_c25, Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_copy3140_c26 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3141_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3141_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w49_32_c26 :  std_logic;
signal bh2587_w50_26_c26 :  std_logic;
signal bh2587_w51_24_c26 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_copy3142_c25, Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_copy3142_c26 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3143_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3143_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w51_25_c26 :  std_logic;
signal bh2587_w52_21_c26 :  std_logic;
signal bh2587_w53_19_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_copy3144_c25, Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_copy3144_c26 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3145_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3145_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w53_20_c26 :  std_logic;
signal bh2587_w54_16_c26 :  std_logic;
signal bh2587_w55_16_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_copy3146_c25, Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_copy3146_c26 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3147_In0_c25 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3147_In1_c25 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_c26 :  std_logic_vector(2 downto 0);
signal bh2587_w55_17_c26 :  std_logic;
signal bh2587_w56_12_c26 :  std_logic;
signal bh2587_w57_12_c26 :  std_logic;
signal Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_copy3148_c25, Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_copy3148_c26 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3149_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3149_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w59_9_c25, bh2587_w59_9_c26 :  std_logic;
signal bh2587_w60_10_c25, bh2587_w60_10_c26 :  std_logic;
signal bh2587_w61_7_c25, bh2587_w61_7_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_copy3150_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3151_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3151_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w61_8_c25, bh2587_w61_8_c26 :  std_logic;
signal bh2587_w62_10_c25, bh2587_w62_10_c26 :  std_logic;
signal bh2587_w63_7_c25, bh2587_w63_7_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_copy3152_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3153_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3153_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w64_11_c25, bh2587_w64_11_c26 :  std_logic;
signal bh2587_w65_7_c25, bh2587_w65_7_c26 :  std_logic;
signal bh2587_w66_11_c25, bh2587_w66_11_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_copy3154_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3155_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3155_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w66_12_c25, bh2587_w66_12_c26 :  std_logic;
signal bh2587_w67_7_c25, bh2587_w67_7_c26 :  std_logic;
signal bh2587_w68_11_c25, bh2587_w68_11_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_copy3156_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3157_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3157_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w68_12_c25, bh2587_w68_12_c26 :  std_logic;
signal bh2587_w69_7_c25, bh2587_w69_7_c26 :  std_logic;
signal bh2587_w70_10_c25, bh2587_w70_10_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_copy3158_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3159_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3159_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w70_11_c25, bh2587_w70_11_c26 :  std_logic;
signal bh2587_w71_6_c25, bh2587_w71_6_c26 :  std_logic;
signal bh2587_w72_10_c25, bh2587_w72_10_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_copy3160_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3161_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3161_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w72_11_c25, bh2587_w72_11_c26 :  std_logic;
signal bh2587_w73_6_c25, bh2587_w73_6_c26 :  std_logic;
signal bh2587_w74_10_c25, bh2587_w74_10_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_copy3162_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3163_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3163_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w74_11_c25, bh2587_w74_11_c26 :  std_logic;
signal bh2587_w75_6_c25, bh2587_w75_6_c26 :  std_logic;
signal bh2587_w76_8_c25, bh2587_w76_8_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_copy3164_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3165_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3165_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w76_9_c25, bh2587_w76_9_c26 :  std_logic;
signal bh2587_w77_4_c25, bh2587_w77_4_c26 :  std_logic;
signal bh2587_w78_6_c25, bh2587_w78_6_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_copy3166_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3167_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3167_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w78_7_c25, bh2587_w78_7_c26 :  std_logic;
signal bh2587_w79_3_c25, bh2587_w79_3_c26 :  std_logic;
signal bh2587_w80_4_c25, bh2587_w80_4_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_copy3168_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3169_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3169_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w80_5_c25, bh2587_w80_5_c26 :  std_logic;
signal bh2587_w81_2_c25, bh2587_w81_2_c26 :  std_logic;
signal bh2587_w82_2_c25, bh2587_w82_2_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_copy3170_c25 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3171_In0_c25 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3171_In1_c25 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_c25 :  std_logic_vector(2 downto 0);
signal bh2587_w82_3_c25, bh2587_w82_3_c26 :  std_logic;
signal bh2587_w83_1_c25, bh2587_w83_1_c26 :  std_logic;
signal bh2587_w84_1_c25, bh2587_w84_1_c26 :  std_logic;
signal Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_copy3172_c25 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh2587_43_c26 :  std_logic_vector(43 downto 0);
signal bitheapFinalAdd_bh2587_In0_c26 :  std_logic_vector(49 downto 0);
signal bitheapFinalAdd_bh2587_In1_c26 :  std_logic_vector(49 downto 0);
signal bitheapFinalAdd_bh2587_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh2587_Out_c26 :  std_logic_vector(49 downto 0);
signal bitheapResult_bh2587_c26 :  std_logic_vector(92 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_21 = '1' then
               bh2587_w39_27_c21 <= bh2587_w39_27_c20;
               bh2587_w40_18_c21 <= bh2587_w40_18_c20;
               bh2587_w41_17_c21 <= bh2587_w41_17_c20;
               bh2587_w42_21_c21 <= bh2587_w42_21_c20;
               bh2587_w43_20_c21 <= bh2587_w43_20_c20;
               bh2587_w44_19_c21 <= bh2587_w44_19_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c20;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c21 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c20;
            end if;
            if ce_22 = '1' then
               bh2587_w39_27_c22 <= bh2587_w39_27_c21;
               bh2587_w40_18_c22 <= bh2587_w40_18_c21;
               bh2587_w41_17_c22 <= bh2587_w41_17_c21;
               bh2587_w42_21_c22 <= bh2587_w42_21_c21;
               bh2587_w43_20_c22 <= bh2587_w43_20_c21;
               bh2587_w44_19_c22 <= bh2587_w44_19_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c21;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c22 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c21;
            end if;
            if ce_23 = '1' then
               bh2587_w39_27_c23 <= bh2587_w39_27_c22;
               bh2587_w40_18_c23 <= bh2587_w40_18_c22;
               bh2587_w41_17_c23 <= bh2587_w41_17_c22;
               bh2587_w42_21_c23 <= bh2587_w42_21_c22;
               bh2587_w43_20_c23 <= bh2587_w43_20_c22;
               bh2587_w44_19_c23 <= bh2587_w44_19_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c22;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c23 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c22;
            end if;
            if ce_24 = '1' then
               bh2587_w39_27_c24 <= bh2587_w39_27_c23;
               bh2587_w40_18_c24 <= bh2587_w40_18_c23;
               bh2587_w41_17_c24 <= bh2587_w41_17_c23;
               bh2587_w42_21_c24 <= bh2587_w42_21_c23;
               bh2587_w43_20_c24 <= bh2587_w43_20_c23;
               bh2587_w44_19_c24 <= bh2587_w44_19_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c23;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c23;
            end if;
            if ce_25 = '1' then
               bh2587_w39_1_c25 <= bh2587_w39_1_c24;
               bh2587_w39_2_c25 <= bh2587_w39_2_c24;
               bh2587_w39_3_c25 <= bh2587_w39_3_c24;
               bh2587_w41_1_c25 <= bh2587_w41_1_c24;
               bh2587_w42_1_c25 <= bh2587_w42_1_c24;
               bh2587_w39_4_c25 <= bh2587_w39_4_c24;
               bh2587_w39_5_c25 <= bh2587_w39_5_c24;
               bh2587_w41_2_c25 <= bh2587_w41_2_c24;
               bh2587_w42_2_c25 <= bh2587_w42_2_c24;
               bh2587_w44_1_c25 <= bh2587_w44_1_c24;
               bh2587_w41_3_c25 <= bh2587_w41_3_c24;
               bh2587_w42_3_c25 <= bh2587_w42_3_c24;
               bh2587_w42_4_c25 <= bh2587_w42_4_c24;
               bh2587_w44_2_c25 <= bh2587_w44_2_c24;
               bh2587_w45_1_c25 <= bh2587_w45_1_c24;
               bh2587_w46_1_c25 <= bh2587_w46_1_c24;
               bh2587_w41_4_c25 <= bh2587_w41_4_c24;
               bh2587_w42_5_c25 <= bh2587_w42_5_c24;
               bh2587_w41_5_c25 <= bh2587_w41_5_c24;
               bh2587_w42_6_c25 <= bh2587_w42_6_c24;
               bh2587_w44_3_c25 <= bh2587_w44_3_c24;
               bh2587_w45_2_c25 <= bh2587_w45_2_c24;
               bh2587_w44_4_c25 <= bh2587_w44_4_c24;
               bh2587_w45_3_c25 <= bh2587_w45_3_c24;
               bh2587_w46_2_c25 <= bh2587_w46_2_c24;
               bh2587_w47_1_c25 <= bh2587_w47_1_c24;
               bh2587_w48_1_c25 <= bh2587_w48_1_c24;
               bh2587_w40_6_c25 <= bh2587_w40_6_c24;
               bh2587_w40_7_c25 <= bh2587_w40_7_c24;
               bh2587_w41_6_c25 <= bh2587_w41_6_c24;
               bh2587_w42_7_c25 <= bh2587_w42_7_c24;
               bh2587_w44_5_c25 <= bh2587_w44_5_c24;
               bh2587_w43_6_c25 <= bh2587_w43_6_c24;
               bh2587_w44_6_c25 <= bh2587_w44_6_c24;
               bh2587_w45_4_c25 <= bh2587_w45_4_c24;
               bh2587_w46_3_c25 <= bh2587_w46_3_c24;
               bh2587_w47_2_c25 <= bh2587_w47_2_c24;
               bh2587_w46_4_c25 <= bh2587_w46_4_c24;
               bh2587_w47_3_c25 <= bh2587_w47_3_c24;
               bh2587_w48_2_c25 <= bh2587_w48_2_c24;
               bh2587_w49_1_c25 <= bh2587_w49_1_c24;
               bh2587_w50_1_c25 <= bh2587_w50_1_c24;
               bh2587_w40_8_c25 <= bh2587_w40_8_c24;
               bh2587_w41_7_c25 <= bh2587_w41_7_c24;
               bh2587_w42_8_c25 <= bh2587_w42_8_c24;
               bh2587_w43_7_c25 <= bh2587_w43_7_c24;
               bh2587_w42_9_c25 <= bh2587_w42_9_c24;
               bh2587_w43_8_c25 <= bh2587_w43_8_c24;
               bh2587_w44_7_c25 <= bh2587_w44_7_c24;
               bh2587_w45_5_c25 <= bh2587_w45_5_c24;
               bh2587_w46_5_c25 <= bh2587_w46_5_c24;
               bh2587_w45_6_c25 <= bh2587_w45_6_c24;
               bh2587_w46_6_c25 <= bh2587_w46_6_c24;
               bh2587_w47_4_c25 <= bh2587_w47_4_c24;
               bh2587_w48_3_c25 <= bh2587_w48_3_c24;
               bh2587_w49_2_c25 <= bh2587_w49_2_c24;
               bh2587_w48_4_c25 <= bh2587_w48_4_c24;
               bh2587_w49_3_c25 <= bh2587_w49_3_c24;
               bh2587_w50_2_c25 <= bh2587_w50_2_c24;
               bh2587_w51_1_c25 <= bh2587_w51_1_c24;
               bh2587_w52_1_c25 <= bh2587_w52_1_c24;
               bh2587_w40_11_c25 <= bh2587_w40_11_c24;
               bh2587_w40_12_c25 <= bh2587_w40_12_c24;
               bh2587_w41_10_c25 <= bh2587_w41_10_c24;
               bh2587_w42_12_c25 <= bh2587_w42_12_c24;
               bh2587_w44_9_c25 <= bh2587_w44_9_c24;
               bh2587_w41_11_c25 <= bh2587_w41_11_c24;
               bh2587_w43_12_c25 <= bh2587_w43_12_c24;
               bh2587_w45_8_c25 <= bh2587_w45_8_c24;
               bh2587_w46_8_c25 <= bh2587_w46_8_c24;
               bh2587_w39_23_c25 <= bh2587_w39_23_c24;
               bh2587_w41_12_c25 <= bh2587_w41_12_c24;
               bh2587_w44_11_c25 <= bh2587_w44_11_c24;
               bh2587_w44_12_c25 <= bh2587_w44_12_c24;
               bh2587_w45_10_c25 <= bh2587_w45_10_c24;
               bh2587_w48_6_c25 <= bh2587_w48_6_c24;
               bh2587_w39_24_c25 <= bh2587_w39_24_c24;
               bh2587_w39_25_c25 <= bh2587_w39_25_c24;
               bh2587_w45_11_c25 <= bh2587_w45_11_c24;
               bh2587_w46_10_c25 <= bh2587_w46_10_c24;
               bh2587_w46_11_c25 <= bh2587_w46_11_c24;
               bh2587_w48_7_c25 <= bh2587_w48_7_c24;
               bh2587_w49_5_c25 <= bh2587_w49_5_c24;
               bh2587_w39_26_c25 <= bh2587_w39_26_c24;
               bh2587_w45_12_c25 <= bh2587_w45_12_c24;
               bh2587_w46_12_c25 <= bh2587_w46_12_c24;
               bh2587_w49_6_c25 <= bh2587_w49_6_c24;
               bh2587_w48_9_c25 <= bh2587_w48_9_c24;
               bh2587_w52_3_c25 <= bh2587_w52_3_c24;
               bh2587_w52_4_c25 <= bh2587_w52_4_c24;
               bh2587_w53_3_c25 <= bh2587_w53_3_c24;
               bh2587_w54_3_c25 <= bh2587_w54_3_c24;
               bh2587_w52_5_c25 <= bh2587_w52_5_c24;
               bh2587_w53_4_c25 <= bh2587_w53_4_c24;
               bh2587_w53_5_c25 <= bh2587_w53_5_c24;
               bh2587_w54_4_c25 <= bh2587_w54_4_c24;
               bh2587_w55_3_c25 <= bh2587_w55_3_c24;
               bh2587_w56_3_c25 <= bh2587_w56_3_c24;
               bh2587_w53_6_c25 <= bh2587_w53_6_c24;
               bh2587_w54_5_c25 <= bh2587_w54_5_c24;
               bh2587_w55_4_c25 <= bh2587_w55_4_c24;
               bh2587_w55_5_c25 <= bh2587_w55_5_c24;
               bh2587_w56_4_c25 <= bh2587_w56_4_c24;
               bh2587_w57_3_c25 <= bh2587_w57_3_c24;
               bh2587_w58_3_c25 <= bh2587_w58_3_c24;
               bh2587_w39_27_c25 <= bh2587_w39_27_c24;
               bh2587_w39_31_c25 <= bh2587_w39_31_c24;
               bh2587_w40_21_c25 <= bh2587_w40_21_c24;
               bh2587_w41_20_c25 <= bh2587_w41_20_c24;
               bh2587_w39_32_c25 <= bh2587_w39_32_c24;
               bh2587_w40_22_c25 <= bh2587_w40_22_c24;
               bh2587_w41_21_c25 <= bh2587_w41_21_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In0_c24;
               bh2587_w40_24_c25 <= bh2587_w40_24_c24;
               bh2587_w41_23_c25 <= bh2587_w41_23_c24;
               bh2587_w42_22_c25 <= bh2587_w42_22_c24;
               bh2587_w40_25_c25 <= bh2587_w40_25_c24;
               bh2587_w41_24_c25 <= bh2587_w41_24_c24;
               bh2587_w42_23_c25 <= bh2587_w42_23_c24;
               bh2587_w41_26_c25 <= bh2587_w41_26_c24;
               bh2587_w42_25_c25 <= bh2587_w42_25_c24;
               bh2587_w43_21_c25 <= bh2587_w43_21_c24;
               bh2587_w42_29_c25 <= bh2587_w42_29_c24;
               bh2587_w43_25_c25 <= bh2587_w43_25_c24;
               bh2587_w44_21_c25 <= bh2587_w44_21_c24;
               bh2587_w42_31_c25 <= bh2587_w42_31_c24;
               bh2587_w43_27_c25 <= bh2587_w43_27_c24;
               bh2587_w43_28_c25 <= bh2587_w43_28_c24;
               bh2587_w44_24_c25 <= bh2587_w44_24_c24;
               bh2587_w45_18_c25 <= bh2587_w45_18_c24;
               bh2587_w43_29_c25 <= bh2587_w43_29_c24;
               bh2587_w45_19_c25 <= bh2587_w45_19_c24;
               bh2587_w43_31_c25 <= bh2587_w43_31_c24;
               bh2587_w45_21_c25 <= bh2587_w45_21_c24;
               bh2587_w45_23_c25 <= bh2587_w45_23_c24;
               bh2587_w46_19_c25 <= bh2587_w46_19_c24;
               bh2587_w45_25_c25 <= bh2587_w45_25_c24;
               bh2587_w46_21_c25 <= bh2587_w46_21_c24;
               bh2587_w47_15_c25 <= bh2587_w47_15_c24;
               bh2587_w46_25_c25 <= bh2587_w46_25_c24;
               bh2587_w47_19_c25 <= bh2587_w47_19_c24;
               bh2587_w48_16_c25 <= bh2587_w48_16_c24;
               bh2587_w47_21_c25 <= bh2587_w47_21_c24;
               bh2587_w48_18_c25 <= bh2587_w48_18_c24;
               bh2587_w49_13_c25 <= bh2587_w49_13_c24;
               Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In0_c24;
               bh2587_w48_21_c25 <= bh2587_w48_21_c24;
               bh2587_w49_16_c25 <= bh2587_w49_16_c24;
               bh2587_w50_11_c25 <= bh2587_w50_11_c24;
               bh2587_w49_19_c25 <= bh2587_w49_19_c24;
               bh2587_w50_14_c25 <= bh2587_w50_14_c24;
               bh2587_w51_10_c25 <= bh2587_w51_10_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In0_c24;
               Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In0_c24;
               bh2587_w51_14_c25 <= bh2587_w51_14_c24;
               bh2587_w52_12_c25 <= bh2587_w52_12_c24;
               bh2587_w53_7_c25 <= bh2587_w53_7_c24;
               bh2587_w52_14_c25 <= bh2587_w52_14_c24;
               bh2587_w53_9_c25 <= bh2587_w53_9_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In0_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In1_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c24;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c24;
            end if;
            if ce_26 = '1' then
               bh2587_w29_0_c26 <= bh2587_w29_0_c25;
               bh2587_w30_0_c26 <= bh2587_w30_0_c25;
               bh2587_w31_0_c26 <= bh2587_w31_0_c25;
               bh2587_w32_0_c26 <= bh2587_w32_0_c25;
               bh2587_w33_0_c26 <= bh2587_w33_0_c25;
               bh2587_w34_0_c26 <= bh2587_w34_0_c25;
               bh2587_w35_0_c26 <= bh2587_w35_0_c25;
               bh2587_w84_0_c26 <= bh2587_w84_0_c25;
               bh2587_w85_0_c26 <= bh2587_w85_0_c25;
               bh2587_w86_0_c26 <= bh2587_w86_0_c25;
               bh2587_w87_0_c26 <= bh2587_w87_0_c25;
               bh2587_w88_0_c26 <= bh2587_w88_0_c25;
               bh2587_w89_0_c26 <= bh2587_w89_0_c25;
               bh2587_w90_0_c26 <= bh2587_w90_0_c25;
               bh2587_w91_0_c26 <= bh2587_w91_0_c25;
               bh2587_w92_0_c26 <= bh2587_w92_0_c25;
               bh2587_w36_2_c26 <= bh2587_w36_2_c25;
               bh2587_w37_3_c26 <= bh2587_w37_3_c25;
               bh2587_w38_5_c26 <= bh2587_w38_5_c25;
               bh2587_w39_36_c26 <= bh2587_w39_36_c25;
               bh2587_w40_32_c26 <= bh2587_w40_32_c25;
               bh2587_w41_36_c26 <= bh2587_w41_36_c25;
               bh2587_w57_11_c26 <= bh2587_w57_11_c25;
               bh2587_w58_12_c26 <= bh2587_w58_12_c25;
               bh2587_w63_6_c26 <= bh2587_w63_6_c25;
               Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_copy3134_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_copy3134_c25;
               Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_copy3136_c26 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_copy3136_c25;
               Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_copy3138_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_copy3138_c25;
               Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_copy3140_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_copy3140_c25;
               Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_copy3142_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_copy3142_c25;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_copy3144_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_copy3144_c25;
               Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_copy3146_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_copy3146_c25;
               Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_copy3148_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_copy3148_c25;
               bh2587_w59_9_c26 <= bh2587_w59_9_c25;
               bh2587_w60_10_c26 <= bh2587_w60_10_c25;
               bh2587_w61_7_c26 <= bh2587_w61_7_c25;
               bh2587_w61_8_c26 <= bh2587_w61_8_c25;
               bh2587_w62_10_c26 <= bh2587_w62_10_c25;
               bh2587_w63_7_c26 <= bh2587_w63_7_c25;
               bh2587_w64_11_c26 <= bh2587_w64_11_c25;
               bh2587_w65_7_c26 <= bh2587_w65_7_c25;
               bh2587_w66_11_c26 <= bh2587_w66_11_c25;
               bh2587_w66_12_c26 <= bh2587_w66_12_c25;
               bh2587_w67_7_c26 <= bh2587_w67_7_c25;
               bh2587_w68_11_c26 <= bh2587_w68_11_c25;
               bh2587_w68_12_c26 <= bh2587_w68_12_c25;
               bh2587_w69_7_c26 <= bh2587_w69_7_c25;
               bh2587_w70_10_c26 <= bh2587_w70_10_c25;
               bh2587_w70_11_c26 <= bh2587_w70_11_c25;
               bh2587_w71_6_c26 <= bh2587_w71_6_c25;
               bh2587_w72_10_c26 <= bh2587_w72_10_c25;
               bh2587_w72_11_c26 <= bh2587_w72_11_c25;
               bh2587_w73_6_c26 <= bh2587_w73_6_c25;
               bh2587_w74_10_c26 <= bh2587_w74_10_c25;
               bh2587_w74_11_c26 <= bh2587_w74_11_c25;
               bh2587_w75_6_c26 <= bh2587_w75_6_c25;
               bh2587_w76_8_c26 <= bh2587_w76_8_c25;
               bh2587_w76_9_c26 <= bh2587_w76_9_c25;
               bh2587_w77_4_c26 <= bh2587_w77_4_c25;
               bh2587_w78_6_c26 <= bh2587_w78_6_c25;
               bh2587_w78_7_c26 <= bh2587_w78_7_c25;
               bh2587_w79_3_c26 <= bh2587_w79_3_c25;
               bh2587_w80_4_c26 <= bh2587_w80_4_c25;
               bh2587_w80_5_c26 <= bh2587_w80_5_c25;
               bh2587_w81_2_c26 <= bh2587_w81_2_c25;
               bh2587_w82_2_c26 <= bh2587_w82_2_c25;
               bh2587_w82_3_c26 <= bh2587_w82_3_c25;
               bh2587_w83_1_c26 <= bh2587_w83_1_c25;
               bh2587_w84_1_c26 <= bh2587_w84_1_c25;
            end if;
         end if;
      end process;
   XX_m2586_c20 <= X ;
   YY_m2586_c24 <= Y ;
   tile_0_X_c20 <= X(45 downto 29);
   tile_0_Y_c24 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid2589
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 X => tile_0_X_c20,
                 Y => tile_0_Y_c24,
                 R => tile_0_output_c25);

   tile_0_filtered_output_c25 <= unsigned(tile_0_output_c25(40 downto 0));
   bh2587_w29_0_c25 <= tile_0_filtered_output_c25(0);
   bh2587_w30_0_c25 <= tile_0_filtered_output_c25(1);
   bh2587_w31_0_c25 <= tile_0_filtered_output_c25(2);
   bh2587_w32_0_c25 <= tile_0_filtered_output_c25(3);
   bh2587_w33_0_c25 <= tile_0_filtered_output_c25(4);
   bh2587_w34_0_c25 <= tile_0_filtered_output_c25(5);
   bh2587_w35_0_c25 <= tile_0_filtered_output_c25(6);
   bh2587_w36_0_c25 <= tile_0_filtered_output_c25(7);
   bh2587_w37_0_c25 <= tile_0_filtered_output_c25(8);
   bh2587_w38_0_c25 <= tile_0_filtered_output_c25(9);
   bh2587_w39_0_c25 <= tile_0_filtered_output_c25(10);
   bh2587_w40_0_c25 <= tile_0_filtered_output_c25(11);
   bh2587_w41_0_c25 <= tile_0_filtered_output_c25(12);
   bh2587_w42_0_c25 <= tile_0_filtered_output_c25(13);
   bh2587_w43_0_c25 <= tile_0_filtered_output_c25(14);
   bh2587_w44_0_c25 <= tile_0_filtered_output_c25(15);
   bh2587_w45_0_c25 <= tile_0_filtered_output_c25(16);
   bh2587_w46_0_c25 <= tile_0_filtered_output_c25(17);
   bh2587_w47_0_c25 <= tile_0_filtered_output_c25(18);
   bh2587_w48_0_c25 <= tile_0_filtered_output_c25(19);
   bh2587_w49_0_c25 <= tile_0_filtered_output_c25(20);
   bh2587_w50_0_c25 <= tile_0_filtered_output_c25(21);
   bh2587_w51_0_c25 <= tile_0_filtered_output_c25(22);
   bh2587_w52_0_c25 <= tile_0_filtered_output_c25(23);
   bh2587_w53_0_c25 <= tile_0_filtered_output_c25(24);
   bh2587_w54_0_c25 <= tile_0_filtered_output_c25(25);
   bh2587_w55_0_c25 <= tile_0_filtered_output_c25(26);
   bh2587_w56_0_c25 <= tile_0_filtered_output_c25(27);
   bh2587_w57_0_c25 <= tile_0_filtered_output_c25(28);
   bh2587_w58_0_c25 <= tile_0_filtered_output_c25(29);
   bh2587_w59_0_c25 <= tile_0_filtered_output_c25(30);
   bh2587_w60_0_c25 <= tile_0_filtered_output_c25(31);
   bh2587_w61_0_c25 <= tile_0_filtered_output_c25(32);
   bh2587_w62_0_c25 <= tile_0_filtered_output_c25(33);
   bh2587_w63_0_c25 <= tile_0_filtered_output_c25(34);
   bh2587_w64_0_c25 <= tile_0_filtered_output_c25(35);
   bh2587_w65_0_c25 <= tile_0_filtered_output_c25(36);
   bh2587_w66_0_c25 <= tile_0_filtered_output_c25(37);
   bh2587_w67_0_c25 <= tile_0_filtered_output_c25(38);
   bh2587_w68_0_c25 <= tile_0_filtered_output_c25(39);
   bh2587_w69_0_c25 <= tile_0_filtered_output_c25(40);
   tile_1_X_c20 <= X(28 downto 28);
   tile_1_Y_c24 <= Y(11 downto 11);
   tile_1_mult: IntMultiplierLUT_1x1_Freq300_uid2591
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_1_X_c20,
                 Y => tile_1_Y_c24,
                 R => tile_1_output_c24);

   tile_1_filtered_output_c24 <= unsigned(tile_1_output_c24(0 downto 0));
   bh2587_w39_1_c24 <= tile_1_filtered_output_c24(0);
   tile_2_X_c20 <= X(26 downto 26);
   tile_2_Y_c24 <= Y(13 downto 13);
   tile_2_mult: IntMultiplierLUT_1x1_Freq300_uid2593
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_2_X_c20,
                 Y => tile_2_Y_c24,
                 R => tile_2_output_c24);

   tile_2_filtered_output_c24 <= unsigned(tile_2_output_c24(0 downto 0));
   bh2587_w39_2_c24 <= tile_2_filtered_output_c24(0);
   tile_3_X_c20 <= X(28 downto 27);
   tile_3_Y_c24 <= Y(13 downto 12);
   tile_3_mult: IntMultiplierLUT_2x2_Freq300_uid2595
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_3_X_c20,
                 Y => tile_3_Y_c24,
                 R => tile_3_output_c24);

   tile_3_filtered_output_c24 <= unsigned(tile_3_output_c24(3 downto 0));
   bh2587_w39_3_c24 <= tile_3_filtered_output_c24(0);
   bh2587_w40_1_c24 <= tile_3_filtered_output_c24(1);
   bh2587_w41_1_c24 <= tile_3_filtered_output_c24(2);
   bh2587_w42_1_c24 <= tile_3_filtered_output_c24(3);
   tile_4_X_c20 <= X(25 downto 25);
   tile_4_Y_c24 <= Y(14 downto 14);
   tile_4_mult: IntMultiplierLUT_1x1_Freq300_uid2600
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_4_X_c20,
                 Y => tile_4_Y_c24,
                 R => tile_4_output_c24);

   tile_4_filtered_output_c24 <= unsigned(tile_4_output_c24(0 downto 0));
   bh2587_w39_4_c24 <= tile_4_filtered_output_c24(0);
   tile_5_X_c20 <= X(25 downto 24);
   tile_5_Y_c24 <= Y(15 downto 15);
   tile_5_mult: IntMultiplierLUT_2x1_Freq300_uid2602
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_5_X_c20,
                 Y => tile_5_Y_c24,
                 R => tile_5_output_c24);

   tile_5_filtered_output_c24 <= unsigned(tile_5_output_c24(1 downto 0));
   bh2587_w39_5_c24 <= tile_5_filtered_output_c24(0);
   bh2587_w40_2_c24 <= tile_5_filtered_output_c24(1);
   tile_6_X_c20 <= X(28 downto 26);
   tile_6_Y_c24 <= Y(15 downto 14);
   tile_6_mult: IntMultiplierLUT_3x2_Freq300_uid2604
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_6_X_c20,
                 Y => tile_6_Y_c24,
                 R => tile_6_output_c24);

   tile_6_filtered_output_c24 <= unsigned(tile_6_output_c24(4 downto 0));
   bh2587_w40_3_c24 <= tile_6_filtered_output_c24(0);
   bh2587_w41_2_c24 <= tile_6_filtered_output_c24(1);
   bh2587_w42_2_c24 <= tile_6_filtered_output_c24(2);
   bh2587_w43_1_c24 <= tile_6_filtered_output_c24(3);
   bh2587_w44_1_c24 <= tile_6_filtered_output_c24(4);
   tile_7_X_c20 <= X(22 downto 22);
   tile_7_Y_c24 <= Y(17 downto 17);
   tile_7_mult: IntMultiplierLUT_1x1_Freq300_uid2609
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_7_X_c20,
                 Y => tile_7_Y_c24,
                 R => tile_7_output_c24);

   tile_7_filtered_output_c24 <= unsigned(tile_7_output_c24(0 downto 0));
   bh2587_w39_6_c24 <= tile_7_filtered_output_c24(0);
   tile_8_X_c20 <= X(25 downto 23);
   tile_8_Y_c24 <= Y(17 downto 16);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid2611
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_8_X_c20,
                 Y => tile_8_Y_c24,
                 R => tile_8_output_c24);

   tile_8_filtered_output_c24 <= unsigned(tile_8_output_c24(4 downto 0));
   bh2587_w39_7_c24 <= tile_8_filtered_output_c24(0);
   bh2587_w40_4_c24 <= tile_8_filtered_output_c24(1);
   bh2587_w41_3_c24 <= tile_8_filtered_output_c24(2);
   bh2587_w42_3_c24 <= tile_8_filtered_output_c24(3);
   bh2587_w43_2_c24 <= tile_8_filtered_output_c24(4);
   tile_9_X_c20 <= X(28 downto 26);
   tile_9_Y_c24 <= Y(17 downto 16);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid2616
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_9_X_c20,
                 Y => tile_9_Y_c24,
                 R => tile_9_output_c24);

   tile_9_filtered_output_c24 <= unsigned(tile_9_output_c24(4 downto 0));
   bh2587_w42_4_c24 <= tile_9_filtered_output_c24(0);
   bh2587_w43_3_c24 <= tile_9_filtered_output_c24(1);
   bh2587_w44_2_c24 <= tile_9_filtered_output_c24(2);
   bh2587_w45_1_c24 <= tile_9_filtered_output_c24(3);
   bh2587_w46_1_c24 <= tile_9_filtered_output_c24(4);
   tile_10_X_c20 <= X(20 downto 20);
   tile_10_Y_c24 <= Y(19 downto 19);
   tile_10_mult: IntMultiplierLUT_1x1_Freq300_uid2621
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_10_X_c20,
                 Y => tile_10_Y_c24,
                 R => tile_10_output_c24);

   tile_10_filtered_output_c24 <= unsigned(tile_10_output_c24(0 downto 0));
   bh2587_w39_8_c24 <= tile_10_filtered_output_c24(0);
   tile_11_X_c20 <= X(22 downto 21);
   tile_11_Y_c24 <= Y(19 downto 18);
   tile_11_mult: IntMultiplierLUT_2x2_Freq300_uid2623
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_11_X_c20,
                 Y => tile_11_Y_c24,
                 R => tile_11_output_c24);

   tile_11_filtered_output_c24 <= unsigned(tile_11_output_c24(3 downto 0));
   bh2587_w39_9_c24 <= tile_11_filtered_output_c24(0);
   bh2587_w40_5_c24 <= tile_11_filtered_output_c24(1);
   bh2587_w41_4_c24 <= tile_11_filtered_output_c24(2);
   bh2587_w42_5_c24 <= tile_11_filtered_output_c24(3);
   tile_12_X_c20 <= X(25 downto 23);
   tile_12_Y_c24 <= Y(19 downto 18);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid2628
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_12_X_c20,
                 Y => tile_12_Y_c24,
                 R => tile_12_output_c24);

   tile_12_filtered_output_c24 <= unsigned(tile_12_output_c24(4 downto 0));
   bh2587_w41_5_c24 <= tile_12_filtered_output_c24(0);
   bh2587_w42_6_c24 <= tile_12_filtered_output_c24(1);
   bh2587_w43_4_c24 <= tile_12_filtered_output_c24(2);
   bh2587_w44_3_c24 <= tile_12_filtered_output_c24(3);
   bh2587_w45_2_c24 <= tile_12_filtered_output_c24(4);
   tile_13_X_c20 <= X(28 downto 26);
   tile_13_Y_c24 <= Y(19 downto 18);
   tile_13_mult: IntMultiplierLUT_3x2_Freq300_uid2633
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_13_X_c20,
                 Y => tile_13_Y_c24,
                 R => tile_13_output_c24);

   tile_13_filtered_output_c24 <= unsigned(tile_13_output_c24(4 downto 0));
   bh2587_w44_4_c24 <= tile_13_filtered_output_c24(0);
   bh2587_w45_3_c24 <= tile_13_filtered_output_c24(1);
   bh2587_w46_2_c24 <= tile_13_filtered_output_c24(2);
   bh2587_w47_1_c24 <= tile_13_filtered_output_c24(3);
   bh2587_w48_1_c24 <= tile_13_filtered_output_c24(4);
   tile_14_X_c20 <= X(19 downto 19);
   tile_14_Y_c24 <= Y(20 downto 20);
   tile_14_mult: IntMultiplierLUT_1x1_Freq300_uid2638
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_14_X_c20,
                 Y => tile_14_Y_c24,
                 R => tile_14_output_c24);

   tile_14_filtered_output_c24 <= unsigned(tile_14_output_c24(0 downto 0));
   bh2587_w39_10_c24 <= tile_14_filtered_output_c24(0);
   tile_15_X_c20 <= X(19 downto 18);
   tile_15_Y_c24 <= Y(21 downto 21);
   tile_15_mult: IntMultiplierLUT_2x1_Freq300_uid2640
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_15_X_c20,
                 Y => tile_15_Y_c24,
                 R => tile_15_output_c24);

   tile_15_filtered_output_c24 <= unsigned(tile_15_output_c24(1 downto 0));
   bh2587_w39_11_c24 <= tile_15_filtered_output_c24(0);
   bh2587_w40_6_c24 <= tile_15_filtered_output_c24(1);
   tile_16_X_c20 <= X(22 downto 20);
   tile_16_Y_c24 <= Y(21 downto 20);
   tile_16_mult: IntMultiplierLUT_3x2_Freq300_uid2642
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_16_X_c20,
                 Y => tile_16_Y_c24,
                 R => tile_16_output_c24);

   tile_16_filtered_output_c24 <= unsigned(tile_16_output_c24(4 downto 0));
   bh2587_w40_7_c24 <= tile_16_filtered_output_c24(0);
   bh2587_w41_6_c24 <= tile_16_filtered_output_c24(1);
   bh2587_w42_7_c24 <= tile_16_filtered_output_c24(2);
   bh2587_w43_5_c24 <= tile_16_filtered_output_c24(3);
   bh2587_w44_5_c24 <= tile_16_filtered_output_c24(4);
   tile_17_X_c20 <= X(25 downto 23);
   tile_17_Y_c24 <= Y(21 downto 20);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid2647
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_17_X_c20,
                 Y => tile_17_Y_c24,
                 R => tile_17_output_c24);

   tile_17_filtered_output_c24 <= unsigned(tile_17_output_c24(4 downto 0));
   bh2587_w43_6_c24 <= tile_17_filtered_output_c24(0);
   bh2587_w44_6_c24 <= tile_17_filtered_output_c24(1);
   bh2587_w45_4_c24 <= tile_17_filtered_output_c24(2);
   bh2587_w46_3_c24 <= tile_17_filtered_output_c24(3);
   bh2587_w47_2_c24 <= tile_17_filtered_output_c24(4);
   tile_18_X_c20 <= X(28 downto 26);
   tile_18_Y_c24 <= Y(21 downto 20);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid2652
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_18_X_c20,
                 Y => tile_18_Y_c24,
                 R => tile_18_output_c24);

   tile_18_filtered_output_c24 <= unsigned(tile_18_output_c24(4 downto 0));
   bh2587_w46_4_c24 <= tile_18_filtered_output_c24(0);
   bh2587_w47_3_c24 <= tile_18_filtered_output_c24(1);
   bh2587_w48_2_c24 <= tile_18_filtered_output_c24(2);
   bh2587_w49_1_c24 <= tile_18_filtered_output_c24(3);
   bh2587_w50_1_c24 <= tile_18_filtered_output_c24(4);
   tile_19_X_c20 <= X(16 downto 16);
   tile_19_Y_c24 <= Y(23 downto 23);
   tile_19_mult: IntMultiplierLUT_1x1_Freq300_uid2657
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_19_X_c20,
                 Y => tile_19_Y_c24,
                 R => tile_19_output_c24);

   tile_19_filtered_output_c24 <= unsigned(tile_19_output_c24(0 downto 0));
   bh2587_w39_12_c24 <= tile_19_filtered_output_c24(0);
   tile_20_X_c20 <= X(19 downto 17);
   tile_20_Y_c24 <= Y(23 downto 22);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid2659
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_20_X_c20,
                 Y => tile_20_Y_c24,
                 R => tile_20_output_c24);

   tile_20_filtered_output_c24 <= unsigned(tile_20_output_c24(4 downto 0));
   bh2587_w39_13_c24 <= tile_20_filtered_output_c24(0);
   bh2587_w40_8_c24 <= tile_20_filtered_output_c24(1);
   bh2587_w41_7_c24 <= tile_20_filtered_output_c24(2);
   bh2587_w42_8_c24 <= tile_20_filtered_output_c24(3);
   bh2587_w43_7_c24 <= tile_20_filtered_output_c24(4);
   tile_21_X_c20 <= X(22 downto 20);
   tile_21_Y_c24 <= Y(23 downto 22);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid2664
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_21_X_c20,
                 Y => tile_21_Y_c24,
                 R => tile_21_output_c24);

   tile_21_filtered_output_c24 <= unsigned(tile_21_output_c24(4 downto 0));
   bh2587_w42_9_c24 <= tile_21_filtered_output_c24(0);
   bh2587_w43_8_c24 <= tile_21_filtered_output_c24(1);
   bh2587_w44_7_c24 <= tile_21_filtered_output_c24(2);
   bh2587_w45_5_c24 <= tile_21_filtered_output_c24(3);
   bh2587_w46_5_c24 <= tile_21_filtered_output_c24(4);
   tile_22_X_c20 <= X(25 downto 23);
   tile_22_Y_c24 <= Y(23 downto 22);
   tile_22_mult: IntMultiplierLUT_3x2_Freq300_uid2669
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_22_X_c20,
                 Y => tile_22_Y_c24,
                 R => tile_22_output_c24);

   tile_22_filtered_output_c24 <= unsigned(tile_22_output_c24(4 downto 0));
   bh2587_w45_6_c24 <= tile_22_filtered_output_c24(0);
   bh2587_w46_6_c24 <= tile_22_filtered_output_c24(1);
   bh2587_w47_4_c24 <= tile_22_filtered_output_c24(2);
   bh2587_w48_3_c24 <= tile_22_filtered_output_c24(3);
   bh2587_w49_2_c24 <= tile_22_filtered_output_c24(4);
   tile_23_X_c20 <= X(28 downto 26);
   tile_23_Y_c24 <= Y(23 downto 22);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid2674
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_23_X_c20,
                 Y => tile_23_Y_c24,
                 R => tile_23_output_c24);

   tile_23_filtered_output_c24 <= unsigned(tile_23_output_c24(4 downto 0));
   bh2587_w48_4_c24 <= tile_23_filtered_output_c24(0);
   bh2587_w49_3_c24 <= tile_23_filtered_output_c24(1);
   bh2587_w50_2_c24 <= tile_23_filtered_output_c24(2);
   bh2587_w51_1_c24 <= tile_23_filtered_output_c24(3);
   bh2587_w52_1_c24 <= tile_23_filtered_output_c24(4);
   tile_24_X_c20 <= X(45 downto 29);
   tile_24_Y_c24 <= Y(46 downto 24);
   tile_24_mult: DSPBlock_17x23_Freq300_uid2679
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 X => tile_24_X_c20,
                 Y => tile_24_Y_c24,
                 R => tile_24_output_c25);

   tile_24_filtered_output_c25 <= unsigned(tile_24_output_c25(39 downto 0));
   bh2587_w53_1_c25 <= tile_24_filtered_output_c25(0);
   bh2587_w54_1_c25 <= tile_24_filtered_output_c25(1);
   bh2587_w55_1_c25 <= tile_24_filtered_output_c25(2);
   bh2587_w56_1_c25 <= tile_24_filtered_output_c25(3);
   bh2587_w57_1_c25 <= tile_24_filtered_output_c25(4);
   bh2587_w58_1_c25 <= tile_24_filtered_output_c25(5);
   bh2587_w59_1_c25 <= tile_24_filtered_output_c25(6);
   bh2587_w60_1_c25 <= tile_24_filtered_output_c25(7);
   bh2587_w61_1_c25 <= tile_24_filtered_output_c25(8);
   bh2587_w62_1_c25 <= tile_24_filtered_output_c25(9);
   bh2587_w63_1_c25 <= tile_24_filtered_output_c25(10);
   bh2587_w64_1_c25 <= tile_24_filtered_output_c25(11);
   bh2587_w65_1_c25 <= tile_24_filtered_output_c25(12);
   bh2587_w66_1_c25 <= tile_24_filtered_output_c25(13);
   bh2587_w67_1_c25 <= tile_24_filtered_output_c25(14);
   bh2587_w68_1_c25 <= tile_24_filtered_output_c25(15);
   bh2587_w69_1_c25 <= tile_24_filtered_output_c25(16);
   bh2587_w70_0_c25 <= tile_24_filtered_output_c25(17);
   bh2587_w71_0_c25 <= tile_24_filtered_output_c25(18);
   bh2587_w72_0_c25 <= tile_24_filtered_output_c25(19);
   bh2587_w73_0_c25 <= tile_24_filtered_output_c25(20);
   bh2587_w74_0_c25 <= tile_24_filtered_output_c25(21);
   bh2587_w75_0_c25 <= tile_24_filtered_output_c25(22);
   bh2587_w76_0_c25 <= tile_24_filtered_output_c25(23);
   bh2587_w77_0_c25 <= tile_24_filtered_output_c25(24);
   bh2587_w78_0_c25 <= tile_24_filtered_output_c25(25);
   bh2587_w79_0_c25 <= tile_24_filtered_output_c25(26);
   bh2587_w80_0_c25 <= tile_24_filtered_output_c25(27);
   bh2587_w81_0_c25 <= tile_24_filtered_output_c25(28);
   bh2587_w82_0_c25 <= tile_24_filtered_output_c25(29);
   bh2587_w83_0_c25 <= tile_24_filtered_output_c25(30);
   bh2587_w84_0_c25 <= tile_24_filtered_output_c25(31);
   bh2587_w85_0_c25 <= tile_24_filtered_output_c25(32);
   bh2587_w86_0_c25 <= tile_24_filtered_output_c25(33);
   bh2587_w87_0_c25 <= tile_24_filtered_output_c25(34);
   bh2587_w88_0_c25 <= tile_24_filtered_output_c25(35);
   bh2587_w89_0_c25 <= tile_24_filtered_output_c25(36);
   bh2587_w90_0_c25 <= tile_24_filtered_output_c25(37);
   bh2587_w91_0_c25 <= tile_24_filtered_output_c25(38);
   bh2587_w92_0_c25 <= tile_24_filtered_output_c25(39);
   tile_25_X_c20 <= X(28 downto 12);
   tile_25_Y_c24 <= Y(46 downto 24);
   tile_25_mult: DSPBlock_17x23_Freq300_uid2681
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 X => tile_25_X_c20,
                 Y => tile_25_Y_c24,
                 R => tile_25_output_c25);

   tile_25_filtered_output_c25 <= unsigned(tile_25_output_c25(39 downto 0));
   bh2587_w36_1_c25 <= tile_25_filtered_output_c25(0);
   bh2587_w37_1_c25 <= tile_25_filtered_output_c25(1);
   bh2587_w38_1_c25 <= tile_25_filtered_output_c25(2);
   bh2587_w39_14_c25 <= tile_25_filtered_output_c25(3);
   bh2587_w40_9_c25 <= tile_25_filtered_output_c25(4);
   bh2587_w41_8_c25 <= tile_25_filtered_output_c25(5);
   bh2587_w42_10_c25 <= tile_25_filtered_output_c25(6);
   bh2587_w43_9_c25 <= tile_25_filtered_output_c25(7);
   bh2587_w44_8_c25 <= tile_25_filtered_output_c25(8);
   bh2587_w45_7_c25 <= tile_25_filtered_output_c25(9);
   bh2587_w46_7_c25 <= tile_25_filtered_output_c25(10);
   bh2587_w47_5_c25 <= tile_25_filtered_output_c25(11);
   bh2587_w48_5_c25 <= tile_25_filtered_output_c25(12);
   bh2587_w49_4_c25 <= tile_25_filtered_output_c25(13);
   bh2587_w50_3_c25 <= tile_25_filtered_output_c25(14);
   bh2587_w51_2_c25 <= tile_25_filtered_output_c25(15);
   bh2587_w52_2_c25 <= tile_25_filtered_output_c25(16);
   bh2587_w53_2_c25 <= tile_25_filtered_output_c25(17);
   bh2587_w54_2_c25 <= tile_25_filtered_output_c25(18);
   bh2587_w55_2_c25 <= tile_25_filtered_output_c25(19);
   bh2587_w56_2_c25 <= tile_25_filtered_output_c25(20);
   bh2587_w57_2_c25 <= tile_25_filtered_output_c25(21);
   bh2587_w58_2_c25 <= tile_25_filtered_output_c25(22);
   bh2587_w59_2_c25 <= tile_25_filtered_output_c25(23);
   bh2587_w60_2_c25 <= tile_25_filtered_output_c25(24);
   bh2587_w61_2_c25 <= tile_25_filtered_output_c25(25);
   bh2587_w62_2_c25 <= tile_25_filtered_output_c25(26);
   bh2587_w63_2_c25 <= tile_25_filtered_output_c25(27);
   bh2587_w64_2_c25 <= tile_25_filtered_output_c25(28);
   bh2587_w65_2_c25 <= tile_25_filtered_output_c25(29);
   bh2587_w66_2_c25 <= tile_25_filtered_output_c25(30);
   bh2587_w67_2_c25 <= tile_25_filtered_output_c25(31);
   bh2587_w68_2_c25 <= tile_25_filtered_output_c25(32);
   bh2587_w69_2_c25 <= tile_25_filtered_output_c25(33);
   bh2587_w70_1_c25 <= tile_25_filtered_output_c25(34);
   bh2587_w71_1_c25 <= tile_25_filtered_output_c25(35);
   bh2587_w72_1_c25 <= tile_25_filtered_output_c25(36);
   bh2587_w73_1_c25 <= tile_25_filtered_output_c25(37);
   bh2587_w74_1_c25 <= tile_25_filtered_output_c25(38);
   bh2587_w75_1_c25 <= tile_25_filtered_output_c25(39);
   tile_26_X_c20 <= X(11 downto 11);
   tile_26_Y_c24 <= Y(28 downto 28);
   tile_26_mult: IntMultiplierLUT_1x1_Freq300_uid2683
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_26_X_c20,
                 Y => tile_26_Y_c24,
                 R => tile_26_output_c24);

   tile_26_filtered_output_c24 <= unsigned(tile_26_output_c24(0 downto 0));
   bh2587_w39_15_c24 <= tile_26_filtered_output_c24(0);
   tile_27_X_c20 <= X(9 downto 9);
   tile_27_Y_c24 <= Y(30 downto 30);
   tile_27_mult: IntMultiplierLUT_1x1_Freq300_uid2685
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_27_X_c20,
                 Y => tile_27_Y_c24,
                 R => tile_27_output_c24);

   tile_27_filtered_output_c24 <= unsigned(tile_27_output_c24(0 downto 0));
   bh2587_w39_16_c24 <= tile_27_filtered_output_c24(0);
   tile_28_X_c20 <= X(11 downto 10);
   tile_28_Y_c24 <= Y(30 downto 29);
   tile_28_mult: IntMultiplierLUT_2x2_Freq300_uid2687
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_28_X_c20,
                 Y => tile_28_Y_c24,
                 R => tile_28_output_c24);

   tile_28_filtered_output_c24 <= unsigned(tile_28_output_c24(3 downto 0));
   bh2587_w39_17_c24 <= tile_28_filtered_output_c24(0);
   bh2587_w40_10_c24 <= tile_28_filtered_output_c24(1);
   bh2587_w41_9_c24 <= tile_28_filtered_output_c24(2);
   bh2587_w42_11_c24 <= tile_28_filtered_output_c24(3);
   tile_29_X_c20 <= X(8 downto 8);
   tile_29_Y_c24 <= Y(31 downto 31);
   tile_29_mult: IntMultiplierLUT_1x1_Freq300_uid2692
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_29_X_c20,
                 Y => tile_29_Y_c24,
                 R => tile_29_output_c24);

   tile_29_filtered_output_c24 <= unsigned(tile_29_output_c24(0 downto 0));
   bh2587_w39_18_c24 <= tile_29_filtered_output_c24(0);
   tile_30_X_c20 <= X(8 downto 7);
   tile_30_Y_c24 <= Y(32 downto 32);
   tile_30_mult: IntMultiplierLUT_2x1_Freq300_uid2694
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_30_X_c20,
                 Y => tile_30_Y_c24,
                 R => tile_30_output_c24);

   tile_30_filtered_output_c24 <= unsigned(tile_30_output_c24(1 downto 0));
   bh2587_w39_19_c24 <= tile_30_filtered_output_c24(0);
   bh2587_w40_11_c24 <= tile_30_filtered_output_c24(1);
   tile_31_X_c20 <= X(11 downto 9);
   tile_31_Y_c24 <= Y(32 downto 31);
   tile_31_mult: IntMultiplierLUT_3x2_Freq300_uid2696
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_31_X_c20,
                 Y => tile_31_Y_c24,
                 R => tile_31_output_c24);

   tile_31_filtered_output_c24 <= unsigned(tile_31_output_c24(4 downto 0));
   bh2587_w40_12_c24 <= tile_31_filtered_output_c24(0);
   bh2587_w41_10_c24 <= tile_31_filtered_output_c24(1);
   bh2587_w42_12_c24 <= tile_31_filtered_output_c24(2);
   bh2587_w43_10_c24 <= tile_31_filtered_output_c24(3);
   bh2587_w44_9_c24 <= tile_31_filtered_output_c24(4);
   tile_32_X_c20 <= X(5 downto 5);
   tile_32_Y_c24 <= Y(34 downto 34);
   tile_32_mult: IntMultiplierLUT_1x1_Freq300_uid2701
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_32_X_c20,
                 Y => tile_32_Y_c24,
                 R => tile_32_output_c24);

   tile_32_filtered_output_c24 <= unsigned(tile_32_output_c24(0 downto 0));
   bh2587_w39_20_c24 <= tile_32_filtered_output_c24(0);
   tile_33_X_c20 <= X(8 downto 6);
   tile_33_Y_c24 <= Y(34 downto 33);
   tile_33_mult: IntMultiplierLUT_3x2_Freq300_uid2703
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_33_X_c20,
                 Y => tile_33_Y_c24,
                 R => tile_33_output_c24);

   tile_33_filtered_output_c24 <= unsigned(tile_33_output_c24(4 downto 0));
   bh2587_w39_21_c24 <= tile_33_filtered_output_c24(0);
   bh2587_w40_13_c24 <= tile_33_filtered_output_c24(1);
   bh2587_w41_11_c24 <= tile_33_filtered_output_c24(2);
   bh2587_w42_13_c24 <= tile_33_filtered_output_c24(3);
   bh2587_w43_11_c24 <= tile_33_filtered_output_c24(4);
   tile_34_X_c20 <= X(11 downto 9);
   tile_34_Y_c24 <= Y(34 downto 33);
   tile_34_mult: IntMultiplierLUT_3x2_Freq300_uid2708
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_34_X_c20,
                 Y => tile_34_Y_c24,
                 R => tile_34_output_c24);

   tile_34_filtered_output_c24 <= unsigned(tile_34_output_c24(4 downto 0));
   bh2587_w42_14_c24 <= tile_34_filtered_output_c24(0);
   bh2587_w43_12_c24 <= tile_34_filtered_output_c24(1);
   bh2587_w44_10_c24 <= tile_34_filtered_output_c24(2);
   bh2587_w45_8_c24 <= tile_34_filtered_output_c24(3);
   bh2587_w46_8_c24 <= tile_34_filtered_output_c24(4);
   tile_35_X_c20 <= X(3 downto 3);
   tile_35_Y_c24 <= Y(36 downto 36);
   tile_35_mult: IntMultiplierLUT_1x1_Freq300_uid2713
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_35_X_c20,
                 Y => tile_35_Y_c24,
                 R => tile_35_output_c24);

   tile_35_filtered_output_c24 <= unsigned(tile_35_output_c24(0 downto 0));
   bh2587_w39_22_c24 <= tile_35_filtered_output_c24(0);
   tile_36_X_c20 <= X(5 downto 4);
   tile_36_Y_c24 <= Y(36 downto 35);
   tile_36_mult: IntMultiplierLUT_2x2_Freq300_uid2715
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_36_X_c20,
                 Y => tile_36_Y_c24,
                 R => tile_36_output_c24);

   tile_36_filtered_output_c24 <= unsigned(tile_36_output_c24(3 downto 0));
   bh2587_w39_23_c24 <= tile_36_filtered_output_c24(0);
   bh2587_w40_14_c24 <= tile_36_filtered_output_c24(1);
   bh2587_w41_12_c24 <= tile_36_filtered_output_c24(2);
   bh2587_w42_15_c24 <= tile_36_filtered_output_c24(3);
   tile_37_X_c20 <= X(8 downto 6);
   tile_37_Y_c24 <= Y(36 downto 35);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid2720
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_37_X_c20,
                 Y => tile_37_Y_c24,
                 R => tile_37_output_c24);

   tile_37_filtered_output_c24 <= unsigned(tile_37_output_c24(4 downto 0));
   bh2587_w41_13_c24 <= tile_37_filtered_output_c24(0);
   bh2587_w42_16_c24 <= tile_37_filtered_output_c24(1);
   bh2587_w43_13_c24 <= tile_37_filtered_output_c24(2);
   bh2587_w44_11_c24 <= tile_37_filtered_output_c24(3);
   bh2587_w45_9_c24 <= tile_37_filtered_output_c24(4);
   tile_38_X_c20 <= X(11 downto 9);
   tile_38_Y_c24 <= Y(36 downto 35);
   tile_38_mult: IntMultiplierLUT_3x2_Freq300_uid2725
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_38_X_c20,
                 Y => tile_38_Y_c24,
                 R => tile_38_output_c24);

   tile_38_filtered_output_c24 <= unsigned(tile_38_output_c24(4 downto 0));
   bh2587_w44_12_c24 <= tile_38_filtered_output_c24(0);
   bh2587_w45_10_c24 <= tile_38_filtered_output_c24(1);
   bh2587_w46_9_c24 <= tile_38_filtered_output_c24(2);
   bh2587_w47_6_c24 <= tile_38_filtered_output_c24(3);
   bh2587_w48_6_c24 <= tile_38_filtered_output_c24(4);
   tile_39_X_c20 <= X(2 downto 2);
   tile_39_Y_c24 <= Y(37 downto 37);
   tile_39_mult: IntMultiplierLUT_1x1_Freq300_uid2730
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_39_X_c20,
                 Y => tile_39_Y_c24,
                 R => tile_39_output_c24);

   tile_39_filtered_output_c24 <= unsigned(tile_39_output_c24(0 downto 0));
   bh2587_w39_24_c24 <= tile_39_filtered_output_c24(0);
   tile_40_X_c20 <= X(2 downto 1);
   tile_40_Y_c24 <= Y(38 downto 38);
   tile_40_mult: IntMultiplierLUT_2x1_Freq300_uid2732
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_40_X_c20,
                 Y => tile_40_Y_c24,
                 R => tile_40_output_c24);

   tile_40_filtered_output_c24 <= unsigned(tile_40_output_c24(1 downto 0));
   bh2587_w39_25_c24 <= tile_40_filtered_output_c24(0);
   bh2587_w40_15_c24 <= tile_40_filtered_output_c24(1);
   tile_41_X_c20 <= X(5 downto 3);
   tile_41_Y_c24 <= Y(38 downto 37);
   tile_41_mult: IntMultiplierLUT_3x2_Freq300_uid2734
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_41_X_c20,
                 Y => tile_41_Y_c24,
                 R => tile_41_output_c24);

   tile_41_filtered_output_c24 <= unsigned(tile_41_output_c24(4 downto 0));
   bh2587_w40_16_c24 <= tile_41_filtered_output_c24(0);
   bh2587_w41_14_c24 <= tile_41_filtered_output_c24(1);
   bh2587_w42_17_c24 <= tile_41_filtered_output_c24(2);
   bh2587_w43_14_c24 <= tile_41_filtered_output_c24(3);
   bh2587_w44_13_c24 <= tile_41_filtered_output_c24(4);
   tile_42_X_c20 <= X(8 downto 6);
   tile_42_Y_c24 <= Y(38 downto 37);
   tile_42_mult: IntMultiplierLUT_3x2_Freq300_uid2739
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_42_X_c20,
                 Y => tile_42_Y_c24,
                 R => tile_42_output_c24);

   tile_42_filtered_output_c24 <= unsigned(tile_42_output_c24(4 downto 0));
   bh2587_w43_15_c24 <= tile_42_filtered_output_c24(0);
   bh2587_w44_14_c24 <= tile_42_filtered_output_c24(1);
   bh2587_w45_11_c24 <= tile_42_filtered_output_c24(2);
   bh2587_w46_10_c24 <= tile_42_filtered_output_c24(3);
   bh2587_w47_7_c24 <= tile_42_filtered_output_c24(4);
   tile_43_X_c20 <= X(11 downto 9);
   tile_43_Y_c24 <= Y(38 downto 37);
   tile_43_mult: IntMultiplierLUT_3x2_Freq300_uid2744
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_43_X_c20,
                 Y => tile_43_Y_c24,
                 R => tile_43_output_c24);

   tile_43_filtered_output_c24 <= unsigned(tile_43_output_c24(4 downto 0));
   bh2587_w46_11_c24 <= tile_43_filtered_output_c24(0);
   bh2587_w47_8_c24 <= tile_43_filtered_output_c24(1);
   bh2587_w48_7_c24 <= tile_43_filtered_output_c24(2);
   bh2587_w49_5_c24 <= tile_43_filtered_output_c24(3);
   bh2587_w50_4_c24 <= tile_43_filtered_output_c24(4);
   tile_44_X_c20 <= X(2 downto 0);
   tile_44_Y_c24 <= Y(40 downto 39);
   tile_44_mult: IntMultiplierLUT_3x2_Freq300_uid2749
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_44_X_c20,
                 Y => tile_44_Y_c24,
                 R => tile_44_output_c24);

   tile_44_filtered_output_c24 <= unsigned(tile_44_output_c24(4 downto 0));
   bh2587_w39_26_c24 <= tile_44_filtered_output_c24(0);
   bh2587_w40_17_c24 <= tile_44_filtered_output_c24(1);
   bh2587_w41_15_c24 <= tile_44_filtered_output_c24(2);
   bh2587_w42_18_c24 <= tile_44_filtered_output_c24(3);
   bh2587_w43_16_c24 <= tile_44_filtered_output_c24(4);
   tile_45_X_c20 <= X(5 downto 3);
   tile_45_Y_c24 <= Y(40 downto 39);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid2754
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_45_X_c20,
                 Y => tile_45_Y_c24,
                 R => tile_45_output_c24);

   tile_45_filtered_output_c24 <= unsigned(tile_45_output_c24(4 downto 0));
   bh2587_w42_19_c24 <= tile_45_filtered_output_c24(0);
   bh2587_w43_17_c24 <= tile_45_filtered_output_c24(1);
   bh2587_w44_15_c24 <= tile_45_filtered_output_c24(2);
   bh2587_w45_12_c24 <= tile_45_filtered_output_c24(3);
   bh2587_w46_12_c24 <= tile_45_filtered_output_c24(4);
   tile_46_X_c20 <= X(8 downto 6);
   tile_46_Y_c24 <= Y(40 downto 39);
   tile_46_mult: IntMultiplierLUT_3x2_Freq300_uid2759
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_46_X_c20,
                 Y => tile_46_Y_c24,
                 R => tile_46_output_c24);

   tile_46_filtered_output_c24 <= unsigned(tile_46_output_c24(4 downto 0));
   bh2587_w45_13_c24 <= tile_46_filtered_output_c24(0);
   bh2587_w46_13_c24 <= tile_46_filtered_output_c24(1);
   bh2587_w47_9_c24 <= tile_46_filtered_output_c24(2);
   bh2587_w48_8_c24 <= tile_46_filtered_output_c24(3);
   bh2587_w49_6_c24 <= tile_46_filtered_output_c24(4);
   tile_47_X_c20 <= X(11 downto 9);
   tile_47_Y_c24 <= Y(40 downto 39);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid2764
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_47_X_c20,
                 Y => tile_47_Y_c24,
                 R => tile_47_output_c24);

   tile_47_filtered_output_c24 <= unsigned(tile_47_output_c24(4 downto 0));
   bh2587_w48_9_c24 <= tile_47_filtered_output_c24(0);
   bh2587_w49_7_c24 <= tile_47_filtered_output_c24(1);
   bh2587_w50_5_c24 <= tile_47_filtered_output_c24(2);
   bh2587_w51_3_c24 <= tile_47_filtered_output_c24(3);
   bh2587_w52_3_c24 <= tile_47_filtered_output_c24(4);
   tile_48_X_c20 <= X(2 downto 0);
   tile_48_Y_c24 <= Y(42 downto 41);
   tile_48_mult: IntMultiplierLUT_3x2_Freq300_uid2769
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_48_X_c20,
                 Y => tile_48_Y_c24,
                 R => tile_48_output_c24);

   tile_48_filtered_output_c24 <= unsigned(tile_48_output_c24(4 downto 0));
   bh2587_w41_16_c24 <= tile_48_filtered_output_c24(0);
   bh2587_w42_20_c24 <= tile_48_filtered_output_c24(1);
   bh2587_w43_18_c24 <= tile_48_filtered_output_c24(2);
   bh2587_w44_16_c24 <= tile_48_filtered_output_c24(3);
   bh2587_w45_14_c24 <= tile_48_filtered_output_c24(4);
   tile_49_X_c20 <= X(5 downto 3);
   tile_49_Y_c24 <= Y(42 downto 41);
   tile_49_mult: IntMultiplierLUT_3x2_Freq300_uid2774
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_49_X_c20,
                 Y => tile_49_Y_c24,
                 R => tile_49_output_c24);

   tile_49_filtered_output_c24 <= unsigned(tile_49_output_c24(4 downto 0));
   bh2587_w44_17_c24 <= tile_49_filtered_output_c24(0);
   bh2587_w45_15_c24 <= tile_49_filtered_output_c24(1);
   bh2587_w46_14_c24 <= tile_49_filtered_output_c24(2);
   bh2587_w47_10_c24 <= tile_49_filtered_output_c24(3);
   bh2587_w48_10_c24 <= tile_49_filtered_output_c24(4);
   tile_50_X_c20 <= X(8 downto 6);
   tile_50_Y_c24 <= Y(42 downto 41);
   tile_50_mult: IntMultiplierLUT_3x2_Freq300_uid2779
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_50_X_c20,
                 Y => tile_50_Y_c24,
                 R => tile_50_output_c24);

   tile_50_filtered_output_c24 <= unsigned(tile_50_output_c24(4 downto 0));
   bh2587_w47_11_c24 <= tile_50_filtered_output_c24(0);
   bh2587_w48_11_c24 <= tile_50_filtered_output_c24(1);
   bh2587_w49_8_c24 <= tile_50_filtered_output_c24(2);
   bh2587_w50_6_c24 <= tile_50_filtered_output_c24(3);
   bh2587_w51_4_c24 <= tile_50_filtered_output_c24(4);
   tile_51_X_c20 <= X(11 downto 9);
   tile_51_Y_c24 <= Y(42 downto 41);
   tile_51_mult: IntMultiplierLUT_3x2_Freq300_uid2784
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_51_X_c20,
                 Y => tile_51_Y_c24,
                 R => tile_51_output_c24);

   tile_51_filtered_output_c24 <= unsigned(tile_51_output_c24(4 downto 0));
   bh2587_w50_7_c24 <= tile_51_filtered_output_c24(0);
   bh2587_w51_5_c24 <= tile_51_filtered_output_c24(1);
   bh2587_w52_4_c24 <= tile_51_filtered_output_c24(2);
   bh2587_w53_3_c24 <= tile_51_filtered_output_c24(3);
   bh2587_w54_3_c24 <= tile_51_filtered_output_c24(4);
   tile_52_X_c20 <= X(2 downto 0);
   tile_52_Y_c24 <= Y(44 downto 43);
   tile_52_mult: IntMultiplierLUT_3x2_Freq300_uid2789
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_52_X_c20,
                 Y => tile_52_Y_c24,
                 R => tile_52_output_c24);

   tile_52_filtered_output_c24 <= unsigned(tile_52_output_c24(4 downto 0));
   bh2587_w43_19_c24 <= tile_52_filtered_output_c24(0);
   bh2587_w44_18_c24 <= tile_52_filtered_output_c24(1);
   bh2587_w45_16_c24 <= tile_52_filtered_output_c24(2);
   bh2587_w46_15_c24 <= tile_52_filtered_output_c24(3);
   bh2587_w47_12_c24 <= tile_52_filtered_output_c24(4);
   tile_53_X_c20 <= X(5 downto 3);
   tile_53_Y_c24 <= Y(44 downto 43);
   tile_53_mult: IntMultiplierLUT_3x2_Freq300_uid2794
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_53_X_c20,
                 Y => tile_53_Y_c24,
                 R => tile_53_output_c24);

   tile_53_filtered_output_c24 <= unsigned(tile_53_output_c24(4 downto 0));
   bh2587_w46_16_c24 <= tile_53_filtered_output_c24(0);
   bh2587_w47_13_c24 <= tile_53_filtered_output_c24(1);
   bh2587_w48_12_c24 <= tile_53_filtered_output_c24(2);
   bh2587_w49_9_c24 <= tile_53_filtered_output_c24(3);
   bh2587_w50_8_c24 <= tile_53_filtered_output_c24(4);
   tile_54_X_c20 <= X(8 downto 6);
   tile_54_Y_c24 <= Y(44 downto 43);
   tile_54_mult: IntMultiplierLUT_3x2_Freq300_uid2799
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_54_X_c20,
                 Y => tile_54_Y_c24,
                 R => tile_54_output_c24);

   tile_54_filtered_output_c24 <= unsigned(tile_54_output_c24(4 downto 0));
   bh2587_w49_10_c24 <= tile_54_filtered_output_c24(0);
   bh2587_w50_9_c24 <= tile_54_filtered_output_c24(1);
   bh2587_w51_6_c24 <= tile_54_filtered_output_c24(2);
   bh2587_w52_5_c24 <= tile_54_filtered_output_c24(3);
   bh2587_w53_4_c24 <= tile_54_filtered_output_c24(4);
   tile_55_X_c20 <= X(11 downto 9);
   tile_55_Y_c24 <= Y(44 downto 43);
   tile_55_mult: IntMultiplierLUT_3x2_Freq300_uid2804
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_55_X_c20,
                 Y => tile_55_Y_c24,
                 R => tile_55_output_c24);

   tile_55_filtered_output_c24 <= unsigned(tile_55_output_c24(4 downto 0));
   bh2587_w52_6_c24 <= tile_55_filtered_output_c24(0);
   bh2587_w53_5_c24 <= tile_55_filtered_output_c24(1);
   bh2587_w54_4_c24 <= tile_55_filtered_output_c24(2);
   bh2587_w55_3_c24 <= tile_55_filtered_output_c24(3);
   bh2587_w56_3_c24 <= tile_55_filtered_output_c24(4);
   tile_56_X_c20 <= X(2 downto 0);
   tile_56_Y_c24 <= Y(46 downto 45);
   tile_56_mult: IntMultiplierLUT_3x2_Freq300_uid2809
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_56_X_c20,
                 Y => tile_56_Y_c24,
                 R => tile_56_output_c24);

   tile_56_filtered_output_c24 <= unsigned(tile_56_output_c24(4 downto 0));
   bh2587_w45_17_c24 <= tile_56_filtered_output_c24(0);
   bh2587_w46_17_c24 <= tile_56_filtered_output_c24(1);
   bh2587_w47_14_c24 <= tile_56_filtered_output_c24(2);
   bh2587_w48_13_c24 <= tile_56_filtered_output_c24(3);
   bh2587_w49_11_c24 <= tile_56_filtered_output_c24(4);
   tile_57_X_c20 <= X(5 downto 3);
   tile_57_Y_c24 <= Y(46 downto 45);
   tile_57_mult: IntMultiplierLUT_3x2_Freq300_uid2814
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_57_X_c20,
                 Y => tile_57_Y_c24,
                 R => tile_57_output_c24);

   tile_57_filtered_output_c24 <= unsigned(tile_57_output_c24(4 downto 0));
   bh2587_w48_14_c24 <= tile_57_filtered_output_c24(0);
   bh2587_w49_12_c24 <= tile_57_filtered_output_c24(1);
   bh2587_w50_10_c24 <= tile_57_filtered_output_c24(2);
   bh2587_w51_7_c24 <= tile_57_filtered_output_c24(3);
   bh2587_w52_7_c24 <= tile_57_filtered_output_c24(4);
   tile_58_X_c20 <= X(8 downto 6);
   tile_58_Y_c24 <= Y(46 downto 45);
   tile_58_mult: IntMultiplierLUT_3x2_Freq300_uid2819
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_58_X_c20,
                 Y => tile_58_Y_c24,
                 R => tile_58_output_c24);

   tile_58_filtered_output_c24 <= unsigned(tile_58_output_c24(4 downto 0));
   bh2587_w51_8_c24 <= tile_58_filtered_output_c24(0);
   bh2587_w52_8_c24 <= tile_58_filtered_output_c24(1);
   bh2587_w53_6_c24 <= tile_58_filtered_output_c24(2);
   bh2587_w54_5_c24 <= tile_58_filtered_output_c24(3);
   bh2587_w55_4_c24 <= tile_58_filtered_output_c24(4);
   tile_59_X_c20 <= X(11 downto 9);
   tile_59_Y_c24 <= Y(46 downto 45);
   tile_59_mult: IntMultiplierLUT_3x2_Freq300_uid2824
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 X => tile_59_X_c20,
                 Y => tile_59_Y_c24,
                 R => tile_59_output_c24);

   tile_59_filtered_output_c24 <= unsigned(tile_59_output_c24(4 downto 0));
   bh2587_w54_6_c24 <= tile_59_filtered_output_c24(0);
   bh2587_w55_5_c24 <= tile_59_filtered_output_c24(1);
   bh2587_w56_4_c24 <= tile_59_filtered_output_c24(2);
   bh2587_w57_3_c24 <= tile_59_filtered_output_c24(3);
   bh2587_w58_3_c24 <= tile_59_filtered_output_c24(4);

   -- Adding the constant bits 
   bh2587_w39_27_c0 <= '1';
   bh2587_w40_18_c0 <= '1';
   bh2587_w41_17_c0 <= '1';
   bh2587_w42_21_c0 <= '1';
   bh2587_w43_20_c0 <= '1';
   bh2587_w44_19_c0 <= '1';


   Compressor_23_3_Freq300_uid2830_bh2587_uid2831_In0_c25 <= "" & bh2587_w36_0_c25 & bh2587_w36_1_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid2831_In1_c25 <= "" & bh2587_w37_0_c25 & bh2587_w37_1_c25;
   bh2587_w36_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_c25(0);
   bh2587_w37_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_c25(1);
   bh2587_w38_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2831: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2831_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2831_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_copy2832_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2831_Out0_copy2832_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid2835_In0_c25 <= "" & bh2587_w38_0_c25 & bh2587_w38_1_c25 & "0";
   bh2587_w38_3_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_c25(0);
   bh2587_w39_28_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid2835: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid2835_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_copy2836_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2835_Out0_copy2836_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2839_In0_c25 <= "" & bh2587_w39_14_c25 & bh2587_w39_27_c25 & bh2587_w39_26_c25 & bh2587_w39_25_c25 & bh2587_w39_24_c25 & bh2587_w39_23_c25;
   bh2587_w39_29_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_c25(0);
   bh2587_w40_19_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_c25(1);
   bh2587_w41_18_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2839: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2839_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_copy2840_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2839_Out0_copy2840_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2841_In0_c25 <= "" & bh2587_w39_0_c25 & bh2587_w39_1_c25 & bh2587_w39_2_c25 & bh2587_w39_3_c25 & bh2587_w39_4_c25 & bh2587_w39_5_c25;
   bh2587_w39_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_c25(0);
   bh2587_w40_20_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_c25(1);
   bh2587_w41_19_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2841: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2841_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_copy2842_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2841_Out0_copy2842_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2843_In0_c24 <= "" & bh2587_w39_22_c24 & bh2587_w39_21_c24 & bh2587_w39_20_c24 & bh2587_w39_19_c24 & bh2587_w39_18_c24 & bh2587_w39_17_c24;
   bh2587_w39_31_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_c24(0);
   bh2587_w40_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_c24(1);
   bh2587_w41_20_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2843: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2843_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_copy2844_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2843_Out0_copy2844_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2845_In0_c24 <= "" & bh2587_w39_6_c24 & bh2587_w39_7_c24 & bh2587_w39_8_c24 & bh2587_w39_9_c24 & bh2587_w39_10_c24 & bh2587_w39_11_c24;
   bh2587_w39_32_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_c24(0);
   bh2587_w40_22_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_c24(1);
   bh2587_w41_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2845: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2845_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_copy2846_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2845_Out0_copy2846_c24; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In0_c24 <= "" & bh2587_w39_15_c24 & bh2587_w39_16_c24 & bh2587_w39_13_c24 & bh2587_w39_12_c24;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In1_c25 <= "" & bh2587_w40_0_c25;
   bh2587_w39_33_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_c25(0);
   bh2587_w40_23_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_c25(1);
   bh2587_w41_22_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2849: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2849_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_copy2850_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2849_Out0_copy2850_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2851_In0_c24 <= "" & bh2587_w40_10_c24 & bh2587_w40_1_c24 & bh2587_w40_2_c24 & bh2587_w40_3_c24 & bh2587_w40_4_c24 & bh2587_w40_5_c24;
   bh2587_w40_24_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_c24(0);
   bh2587_w41_23_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_c24(1);
   bh2587_w42_22_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2851: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2851_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_copy2852_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2851_Out0_copy2852_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2853_In0_c24 <= "" & bh2587_w40_18_c24 & bh2587_w40_17_c24 & bh2587_w40_16_c24 & bh2587_w40_15_c24 & bh2587_w40_14_c24 & bh2587_w40_13_c24;
   bh2587_w40_25_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_c24(0);
   bh2587_w41_24_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_c24(1);
   bh2587_w42_23_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2853: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2853_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_copy2854_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2853_Out0_copy2854_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2855_In0_c25 <= "" & bh2587_w40_6_c25 & bh2587_w40_7_c25 & bh2587_w40_8_c25 & bh2587_w40_9_c25 & bh2587_w40_11_c25 & bh2587_w40_12_c25;
   bh2587_w40_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_c25(0);
   bh2587_w41_25_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_c25(1);
   bh2587_w42_24_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2855: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2855_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_copy2856_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2855_Out0_copy2856_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2857_In0_c24 <= "" & bh2587_w41_9_c24 & bh2587_w41_17_c24 & bh2587_w41_16_c24 & bh2587_w41_15_c24 & bh2587_w41_14_c24 & bh2587_w41_13_c24;
   bh2587_w41_26_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_c24(0);
   bh2587_w42_25_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_c24(1);
   bh2587_w43_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2857: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2857_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_copy2858_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2857_Out0_copy2858_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2859_In0_c25 <= "" & bh2587_w41_0_c25 & bh2587_w41_1_c25 & bh2587_w41_2_c25 & bh2587_w41_3_c25 & bh2587_w41_4_c25 & bh2587_w41_5_c25;
   bh2587_w41_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_c25(0);
   bh2587_w42_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_c25(1);
   bh2587_w43_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2859: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2859_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_copy2860_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2859_Out0_copy2860_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2861_In0_c25 <= "" & bh2587_w41_12_c25 & bh2587_w41_11_c25 & bh2587_w41_10_c25 & bh2587_w41_8_c25 & bh2587_w41_7_c25 & bh2587_w41_6_c25;
   bh2587_w41_28_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_c25(0);
   bh2587_w42_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_c25(1);
   bh2587_w43_23_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2861: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2861_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_copy2862_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2861_Out0_copy2862_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2863_In0_c25 <= "" & bh2587_w42_0_c25 & bh2587_w42_1_c25 & bh2587_w42_2_c25 & bh2587_w42_3_c25 & bh2587_w42_4_c25 & bh2587_w42_5_c25;
   bh2587_w42_28_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_c25(0);
   bh2587_w43_24_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_c25(1);
   bh2587_w44_20_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2863: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2863_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_copy2864_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2863_Out0_copy2864_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2865_In0_c24 <= "" & bh2587_w42_11_c24 & bh2587_w42_21_c24 & bh2587_w42_20_c24 & bh2587_w42_19_c24 & bh2587_w42_18_c24 & bh2587_w42_17_c24;
   bh2587_w42_29_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_c24(0);
   bh2587_w43_25_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_c24(1);
   bh2587_w44_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2865: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2865_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_copy2866_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2865_Out0_copy2866_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2867_In0_c25 <= "" & bh2587_w42_6_c25 & bh2587_w42_7_c25 & bh2587_w42_8_c25 & bh2587_w42_9_c25 & bh2587_w42_10_c25 & bh2587_w42_12_c25;
   bh2587_w42_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_c25(0);
   bh2587_w43_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_c25(1);
   bh2587_w44_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2867: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2867_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_copy2868_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2867_Out0_copy2868_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In0_c24 <= "" & bh2587_w42_16_c24 & bh2587_w42_15_c24 & bh2587_w42_14_c24 & bh2587_w42_13_c24;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c0 <= "" & "0";
   bh2587_w42_31_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_c24(0);
   bh2587_w43_27_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_c24(1);
   bh2587_w44_23_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_c24(2);
   Compressor_14_3_Freq300_uid2848_uid2869: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In0_c24,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2869_In1_c24,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_copy2870_c24);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_c24 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2869_Out0_copy2870_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2871_In0_c24 <= "" & bh2587_w43_10_c24 & bh2587_w43_1_c24 & bh2587_w43_2_c24 & bh2587_w43_3_c24 & bh2587_w43_4_c24 & bh2587_w43_5_c24;
   bh2587_w43_28_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_c24(0);
   bh2587_w44_24_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_c24(1);
   bh2587_w45_18_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2871: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2871_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_copy2872_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2871_Out0_copy2872_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2873_In0_c24 <= "" & bh2587_w43_11_c24 & bh2587_w43_20_c24 & bh2587_w43_19_c24 & bh2587_w43_18_c24 & bh2587_w43_17_c24 & bh2587_w43_16_c24;
   bh2587_w43_29_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_c24(0);
   bh2587_w44_25_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_c24(1);
   bh2587_w45_19_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2873: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2873_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_copy2874_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2873_Out0_copy2874_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2875_In0_c25 <= "" & bh2587_w43_6_c25 & bh2587_w43_7_c25 & bh2587_w43_8_c25 & bh2587_w43_9_c25 & bh2587_w43_0_c25 & bh2587_w43_12_c25;
   bh2587_w43_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_c25(0);
   bh2587_w44_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_c25(1);
   bh2587_w45_20_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2875: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2875_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_copy2876_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2875_Out0_copy2876_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2877_In0_c24 <= "" & bh2587_w43_15_c24 & bh2587_w43_14_c24 & bh2587_w43_13_c24;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2877_In1_c24 <= "" & bh2587_w44_10_c24 & bh2587_w44_19_c24;
   bh2587_w43_31_c24 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_c24(0);
   bh2587_w44_27_c24 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_c24(1);
   bh2587_w45_21_c24 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_c24(2);
   Compressor_23_3_Freq300_uid2830_uid2877: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2877_In0_c24,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2877_In1_c24,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_copy2878_c24);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_c24 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2877_Out0_copy2878_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2879_In0_c25 <= "" & bh2587_w44_0_c25 & bh2587_w44_1_c25 & bh2587_w44_2_c25 & bh2587_w44_3_c25 & bh2587_w44_4_c25 & bh2587_w44_5_c25;
   bh2587_w44_28_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_c25(0);
   bh2587_w45_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_c25(1);
   bh2587_w46_18_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2879: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2879_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_copy2880_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2879_Out0_copy2880_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2881_In0_c24 <= "" & bh2587_w44_18_c24 & bh2587_w44_17_c24 & bh2587_w44_16_c24 & bh2587_w44_15_c24 & bh2587_w44_14_c24 & bh2587_w44_13_c24;
   bh2587_w44_29_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_c24(0);
   bh2587_w45_23_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_c24(1);
   bh2587_w46_19_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2881: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2881_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_copy2882_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2881_Out0_copy2882_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2883_In0_c25 <= "" & bh2587_w44_6_c25 & bh2587_w44_7_c25 & bh2587_w44_8_c25 & bh2587_w44_9_c25 & bh2587_w44_11_c25 & bh2587_w44_12_c25;
   bh2587_w44_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_c25(0);
   bh2587_w45_24_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_c25(1);
   bh2587_w46_20_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2883: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2883_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_copy2884_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2883_Out0_copy2884_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2885_In0_c24 <= "" & bh2587_w45_9_c24 & bh2587_w45_17_c24 & bh2587_w45_16_c24 & bh2587_w45_15_c24 & bh2587_w45_14_c24 & bh2587_w45_13_c24;
   bh2587_w45_25_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_c24(0);
   bh2587_w46_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_c24(1);
   bh2587_w47_15_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2885: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2885_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_copy2886_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2885_Out0_copy2886_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2887_In0_c25 <= "" & bh2587_w45_0_c25 & bh2587_w45_1_c25 & bh2587_w45_2_c25 & bh2587_w45_3_c25 & bh2587_w45_4_c25 & bh2587_w45_5_c25;
   bh2587_w45_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_c25(0);
   bh2587_w46_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_c25(1);
   bh2587_w47_16_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2887: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2887_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_copy2888_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2887_Out0_copy2888_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2889_In0_c25 <= "" & bh2587_w45_12_c25 & bh2587_w45_11_c25 & bh2587_w45_10_c25 & bh2587_w45_8_c25 & bh2587_w45_7_c25 & bh2587_w45_6_c25;
   bh2587_w45_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_c25(0);
   bh2587_w46_23_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_c25(1);
   bh2587_w47_17_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2889: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2889_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_copy2890_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2889_Out0_copy2890_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2891_In0_c25 <= "" & bh2587_w46_0_c25 & bh2587_w46_1_c25 & bh2587_w46_2_c25 & bh2587_w46_3_c25 & bh2587_w46_4_c25 & bh2587_w46_5_c25;
   bh2587_w46_24_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_c25(0);
   bh2587_w47_18_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_c25(1);
   bh2587_w48_15_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2891: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2891_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_copy2892_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2891_Out0_copy2892_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2893_In0_c24 <= "" & bh2587_w46_9_c24 & bh2587_w46_17_c24 & bh2587_w46_16_c24 & bh2587_w46_15_c24 & bh2587_w46_14_c24 & bh2587_w46_13_c24;
   bh2587_w46_25_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_c24(0);
   bh2587_w47_19_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_c24(1);
   bh2587_w48_16_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2893: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2893_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_copy2894_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2893_Out0_copy2894_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2895_In0_c25 <= "" & bh2587_w46_6_c25 & bh2587_w46_7_c25 & bh2587_w46_8_c25 & bh2587_w46_10_c25 & bh2587_w46_11_c25 & bh2587_w46_12_c25;
   bh2587_w46_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_c25(0);
   bh2587_w47_20_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_c25(1);
   bh2587_w48_17_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2895: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2895_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_copy2896_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2895_Out0_copy2896_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2897_In0_c24 <= "" & bh2587_w47_8_c24 & bh2587_w47_14_c24 & bh2587_w47_13_c24 & bh2587_w47_12_c24 & bh2587_w47_11_c24 & bh2587_w47_10_c24;
   bh2587_w47_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_c24(0);
   bh2587_w48_18_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_c24(1);
   bh2587_w49_13_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2897: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2897_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_copy2898_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2897_Out0_copy2898_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2899_In0_c25 <= "" & bh2587_w47_0_c25 & bh2587_w47_1_c25 & bh2587_w47_2_c25 & bh2587_w47_3_c25 & bh2587_w47_4_c25 & bh2587_w47_5_c25;
   bh2587_w47_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_c25(0);
   bh2587_w48_19_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_c25(1);
   bh2587_w49_14_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2899: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2899_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_copy2900_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2899_Out0_copy2900_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In0_c24 <= "" & bh2587_w47_9_c24 & bh2587_w47_7_c24 & bh2587_w47_6_c24;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In1_c25 <= "" & bh2587_w48_0_c25 & bh2587_w48_1_c25;
   bh2587_w47_23_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_c25(0);
   bh2587_w48_20_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_c25(1);
   bh2587_w49_15_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2901: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2901_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_copy2902_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2901_Out0_copy2902_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2903_In0_c24 <= "" & bh2587_w48_8_c24 & bh2587_w48_14_c24 & bh2587_w48_13_c24 & bh2587_w48_12_c24 & bh2587_w48_11_c24 & bh2587_w48_10_c24;
   bh2587_w48_21_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_c24(0);
   bh2587_w49_16_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_c24(1);
   bh2587_w50_11_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2903: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2903_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_copy2904_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2903_Out0_copy2904_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2905_In0_c25 <= "" & bh2587_w48_2_c25 & bh2587_w48_3_c25 & bh2587_w48_4_c25 & bh2587_w48_5_c25 & bh2587_w48_6_c25 & bh2587_w48_7_c25;
   bh2587_w48_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_c25(0);
   bh2587_w49_17_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_c25(1);
   bh2587_w50_12_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2905: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2905_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_copy2906_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2905_Out0_copy2906_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2907_In0_c25 <= "" & bh2587_w49_0_c25 & bh2587_w49_1_c25 & bh2587_w49_2_c25 & bh2587_w49_3_c25 & bh2587_w49_4_c25 & bh2587_w49_5_c25;
   bh2587_w49_18_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_c25(0);
   bh2587_w50_13_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_c25(1);
   bh2587_w51_9_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2907: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2907_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_copy2908_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2907_Out0_copy2908_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2909_In0_c24 <= "" & bh2587_w49_8_c24 & bh2587_w49_12_c24 & bh2587_w49_11_c24 & bh2587_w49_10_c24 & bh2587_w49_9_c24 & bh2587_w49_7_c24;
   bh2587_w49_19_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_c24(0);
   bh2587_w50_14_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_c24(1);
   bh2587_w51_10_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2909: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2909_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_copy2910_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2909_Out0_copy2910_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2911_In0_c25 <= "" & bh2587_w50_0_c25 & bh2587_w50_1_c25 & bh2587_w50_2_c25 & bh2587_w50_3_c25 & "0" & "0";
   bh2587_w50_15_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_c25(0);
   bh2587_w51_11_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_c25(1);
   bh2587_w52_9_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2911: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2911_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_copy2912_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2911_Out0_copy2912_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In0_c24 <= "" & bh2587_w50_4_c24 & bh2587_w50_5_c24 & bh2587_w50_6_c24 & bh2587_w50_7_c24;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In1_c25 <= "" & bh2587_w51_0_c25;
   bh2587_w50_16_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_c25(0);
   bh2587_w51_12_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_c25(1);
   bh2587_w52_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2913: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2913_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_copy2914_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2913_Out0_copy2914_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In0_c24 <= "" & bh2587_w50_8_c24 & bh2587_w50_10_c24 & bh2587_w50_9_c24;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In1_c25 <= "" & bh2587_w51_1_c25 & bh2587_w51_2_c25;
   bh2587_w50_17_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_c25(0);
   bh2587_w51_13_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_c25(1);
   bh2587_w52_11_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2915: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2915_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_copy2916_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2915_Out0_copy2916_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2917_In0_c24 <= "" & bh2587_w51_3_c24 & bh2587_w51_4_c24 & bh2587_w51_5_c24 & bh2587_w51_6_c24 & bh2587_w51_7_c24 & bh2587_w51_8_c24;
   bh2587_w51_14_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_c24(0);
   bh2587_w52_12_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_c24(1);
   bh2587_w53_7_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_c24(2);
   Compressor_6_3_Freq300_uid2838_uid2917: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2917_In0_c24,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_copy2918_c24);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_c24 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2917_Out0_copy2918_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2919_In0_c25 <= "" & bh2587_w52_0_c25 & bh2587_w52_1_c25 & bh2587_w52_2_c25 & bh2587_w52_3_c25 & bh2587_w52_4_c25 & bh2587_w52_5_c25;
   bh2587_w52_13_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_c25(0);
   bh2587_w53_8_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_c25(1);
   bh2587_w54_7_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2919: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2919_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_copy2920_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2919_Out0_copy2920_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid2921_In0_c24 <= "" & bh2587_w52_6_c24 & bh2587_w52_7_c24 & bh2587_w52_8_c24;
   bh2587_w52_14_c24 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_c24(0);
   bh2587_w53_9_c24 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_c24(1);
   Compressor_3_2_Freq300_uid2834_uid2921: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid2921_In0_c24,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_copy2922_c24);
   Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_c24 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2921_Out0_copy2922_c24; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2923_In0_c25 <= "" & bh2587_w53_0_c25 & bh2587_w53_1_c25 & bh2587_w53_2_c25 & bh2587_w53_3_c25 & bh2587_w53_4_c25 & bh2587_w53_5_c25;
   bh2587_w53_10_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_c25(0);
   bh2587_w54_8_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_c25(1);
   bh2587_w55_6_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2923: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2923_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_copy2924_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2923_Out0_copy2924_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2925_In0_c25 <= "" & bh2587_w54_0_c25 & bh2587_w54_1_c25 & bh2587_w54_2_c25 & bh2587_w54_3_c25 & bh2587_w54_4_c25 & bh2587_w54_5_c25;
   bh2587_w54_9_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_c25(0);
   bh2587_w55_7_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_c25(1);
   bh2587_w56_5_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2925: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2925_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_copy2926_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2925_Out0_copy2926_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2927_In0_c25 <= "" & bh2587_w55_0_c25 & bh2587_w55_1_c25 & bh2587_w55_2_c25 & bh2587_w55_3_c25 & bh2587_w55_4_c25 & bh2587_w55_5_c25;
   bh2587_w55_8_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_c25(0);
   bh2587_w56_6_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_c25(1);
   bh2587_w57_4_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2927: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2927_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_copy2928_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2927_Out0_copy2928_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2929_In0_c25 <= "" & bh2587_w56_0_c25 & bh2587_w56_1_c25 & bh2587_w56_2_c25 & bh2587_w56_3_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2929_In1_c25 <= "" & bh2587_w57_0_c25;
   bh2587_w56_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_c25(0);
   bh2587_w57_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_c25(1);
   bh2587_w58_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2929: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2929_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2929_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_copy2930_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2929_Out0_copy2930_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid2931_In0_c25 <= "" & bh2587_w57_1_c25 & bh2587_w57_2_c25 & bh2587_w57_3_c25;
   bh2587_w57_6_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_c25(0);
   bh2587_w58_5_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid2931: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid2931_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_copy2932_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2931_Out0_copy2932_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In0_c25 <= "" & bh2587_w58_0_c25 & bh2587_w58_1_c25 & bh2587_w58_2_c25 & bh2587_w58_3_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c0 <= "" & "0";
   bh2587_w58_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_c25(0);
   bh2587_w59_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_c25(1);
   bh2587_w60_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2933: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2933_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_copy2934_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2933_Out0_copy2934_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid2935_In0_c25 <= "" & bh2587_w59_0_c25 & bh2587_w59_1_c25 & bh2587_w59_2_c25;
   bh2587_w59_4_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_c25(0);
   bh2587_w60_4_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid2935: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid2935_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_copy2936_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2935_Out0_copy2936_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2937_In0_c25 <= "" & bh2587_w60_0_c25 & bh2587_w60_1_c25 & bh2587_w60_2_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2937_In1_c25 <= "" & bh2587_w61_0_c25 & bh2587_w61_1_c25;
   bh2587_w60_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_c25(0);
   bh2587_w61_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_c25(1);
   bh2587_w62_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2937: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2937_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2937_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_copy2938_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2937_Out0_copy2938_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2939_In0_c25 <= "" & bh2587_w62_0_c25 & bh2587_w62_1_c25 & bh2587_w62_2_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2939_In1_c25 <= "" & bh2587_w63_0_c25 & bh2587_w63_1_c25;
   bh2587_w62_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_c25(0);
   bh2587_w63_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_c25(1);
   bh2587_w64_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2939: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2939_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2939_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_copy2940_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2939_Out0_copy2940_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2941_In0_c25 <= "" & bh2587_w64_0_c25 & bh2587_w64_1_c25 & bh2587_w64_2_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2941_In1_c25 <= "" & bh2587_w65_0_c25 & bh2587_w65_1_c25;
   bh2587_w64_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_c25(0);
   bh2587_w65_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_c25(1);
   bh2587_w66_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2941: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2941_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2941_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_copy2942_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2941_Out0_copy2942_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2943_In0_c25 <= "" & bh2587_w66_0_c25 & bh2587_w66_1_c25 & bh2587_w66_2_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2943_In1_c25 <= "" & bh2587_w67_0_c25 & bh2587_w67_1_c25;
   bh2587_w66_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_c25(0);
   bh2587_w67_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_c25(1);
   bh2587_w68_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2943: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2943_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2943_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_copy2944_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2943_Out0_copy2944_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2945_In0_c25 <= "" & bh2587_w68_0_c25 & bh2587_w68_1_c25 & bh2587_w68_2_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2945_In1_c25 <= "" & bh2587_w69_0_c25 & bh2587_w69_1_c25;
   bh2587_w68_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_c25(0);
   bh2587_w69_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_c25(1);
   bh2587_w70_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2945: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2945_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2945_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_copy2946_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2945_Out0_copy2946_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2947_In0_c25 <= "" & bh2587_w70_0_c25 & bh2587_w70_1_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid2947_In1_c25 <= "" & bh2587_w71_0_c25 & bh2587_w71_1_c25;
   bh2587_w70_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_c25(0);
   bh2587_w71_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_c25(1);
   bh2587_w72_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2947: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2947_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2947_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_copy2948_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2947_Out0_copy2948_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2949_In0_c25 <= "" & bh2587_w72_0_c25 & bh2587_w72_1_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid2949_In1_c25 <= "" & bh2587_w73_0_c25 & bh2587_w73_1_c25;
   bh2587_w72_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_c25(0);
   bh2587_w73_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_c25(1);
   bh2587_w74_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2949: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2949_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2949_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_copy2950_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2949_Out0_copy2950_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2951_In0_c25 <= "" & bh2587_w74_0_c25 & bh2587_w74_1_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid2951_In1_c25 <= "" & bh2587_w75_0_c25 & bh2587_w75_1_c25;
   bh2587_w74_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_c25(0);
   bh2587_w75_2_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_c25(1);
   bh2587_w76_1_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2951: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2951_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2951_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_copy2952_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2951_Out0_copy2952_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2953_In0_c25 <= "" & bh2587_w37_2_c25 & "0" & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid2953_In1_c25 <= "" & bh2587_w38_2_c25 & bh2587_w38_3_c25;
   bh2587_w37_3_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_c25(0);
   bh2587_w38_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_c25(1);
   bh2587_w39_34_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2953: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2953_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2953_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_copy2954_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2953_Out0_copy2954_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2955_In0_c25 <= "" & bh2587_w39_28_c25 & bh2587_w39_30_c25 & bh2587_w39_32_c25 & bh2587_w39_29_c25 & bh2587_w39_31_c25 & bh2587_w39_33_c25;
   bh2587_w39_35_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_c25(0);
   bh2587_w40_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_c25(1);
   bh2587_w41_29_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2955: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2955_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_copy2956_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2955_Out0_copy2956_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2957_In0_c25 <= "" & bh2587_w40_26_c25 & bh2587_w40_24_c25 & bh2587_w40_22_c25 & bh2587_w40_20_c25 & "0" & "0";
   bh2587_w40_28_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_c25(0);
   bh2587_w41_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_c25(1);
   bh2587_w42_32_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2957: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2957_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_copy2958_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2957_Out0_copy2958_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2959_In0_c25 <= "" & bh2587_w40_19_c25 & bh2587_w40_21_c25 & bh2587_w40_23_c25 & bh2587_w40_25_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2959_In1_c25 <= "" & bh2587_w41_27_c25;
   bh2587_w40_29_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_c25(0);
   bh2587_w41_31_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_c25(1);
   bh2587_w42_33_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2959: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2959_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2959_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_copy2960_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2959_Out0_copy2960_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2961_In0_c25 <= "" & bh2587_w41_25_c25 & bh2587_w41_23_c25 & bh2587_w41_21_c25 & bh2587_w41_19_c25 & bh2587_w41_18_c25 & bh2587_w41_20_c25;
   bh2587_w41_32_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_c25(0);
   bh2587_w42_34_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_c25(1);
   bh2587_w43_32_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2961: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2961_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_copy2962_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2961_Out0_copy2962_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2963_In0_c25 <= "" & bh2587_w41_22_c25 & bh2587_w41_24_c25 & bh2587_w41_26_c25 & bh2587_w41_28_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2963_In1_c25 <= "" & bh2587_w42_30_c25;
   bh2587_w41_33_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_c25(0);
   bh2587_w42_35_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_c25(1);
   bh2587_w43_33_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2963: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2963_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2963_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_copy2964_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2963_Out0_copy2964_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2965_In0_c25 <= "" & bh2587_w42_28_c25 & bh2587_w42_26_c25 & bh2587_w42_24_c25 & bh2587_w42_22_c25 & bh2587_w42_23_c25 & bh2587_w42_25_c25;
   bh2587_w42_36_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_c25(0);
   bh2587_w43_34_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_c25(1);
   bh2587_w44_31_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2965: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2965_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_copy2966_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2965_Out0_copy2966_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid2967_In0_c25 <= "" & bh2587_w42_27_c25 & bh2587_w42_29_c25 & bh2587_w42_31_c25;
   bh2587_w42_37_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_c25(0);
   bh2587_w43_35_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid2967: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid2967_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_copy2968_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid2967_Out0_copy2968_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2969_In0_c25 <= "" & bh2587_w43_30_c25 & bh2587_w43_28_c25 & bh2587_w43_26_c25 & bh2587_w43_24_c25 & bh2587_w43_22_c25 & bh2587_w43_21_c25;
   bh2587_w43_36_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_c25(0);
   bh2587_w44_32_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_c25(1);
   bh2587_w45_28_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2969: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2969_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_copy2970_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2969_Out0_copy2970_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2971_In0_c25 <= "" & bh2587_w43_23_c25 & bh2587_w43_25_c25 & bh2587_w43_27_c25 & bh2587_w43_29_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2971_In1_c25 <= "" & bh2587_w44_30_c25;
   bh2587_w43_37_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_c25(0);
   bh2587_w44_33_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_c25(1);
   bh2587_w45_29_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2971: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2971_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2971_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_copy2972_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2971_Out0_copy2972_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2973_In0_c25 <= "" & bh2587_w44_28_c25 & bh2587_w44_26_c25 & bh2587_w44_24_c25 & bh2587_w44_22_c25 & bh2587_w44_20_c25 & bh2587_w44_21_c25;
   bh2587_w44_34_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_c25(0);
   bh2587_w45_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_c25(1);
   bh2587_w46_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2973: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2973_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_copy2974_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2973_Out0_copy2974_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In0_c24 <= "" & bh2587_w44_23_c24 & bh2587_w44_25_c24 & bh2587_w44_27_c24 & bh2587_w44_29_c24;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In1_c25 <= "" & bh2587_w45_26_c25;
   bh2587_w44_35_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_c25(0);
   bh2587_w45_31_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_c25(1);
   bh2587_w46_28_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2975: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2975_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_copy2976_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2975_Out0_copy2976_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2977_In0_c25 <= "" & bh2587_w45_24_c25 & bh2587_w45_22_c25 & bh2587_w45_20_c25 & bh2587_w45_18_c25 & bh2587_w45_19_c25 & bh2587_w45_21_c25;
   bh2587_w45_32_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_c25(0);
   bh2587_w46_29_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_c25(1);
   bh2587_w47_24_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2977: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2977_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_copy2978_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2977_Out0_copy2978_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2979_In0_c25 <= "" & bh2587_w45_23_c25 & bh2587_w45_25_c25 & bh2587_w45_27_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2979_In1_c25 <= "" & bh2587_w46_26_c25 & bh2587_w46_24_c25;
   bh2587_w45_33_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_c25(0);
   bh2587_w46_30_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_c25(1);
   bh2587_w47_25_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2979: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2979_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2979_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_copy2980_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2979_Out0_copy2980_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2981_In0_c25 <= "" & bh2587_w46_22_c25 & bh2587_w46_20_c25 & bh2587_w46_18_c25 & bh2587_w46_19_c25 & bh2587_w46_21_c25 & bh2587_w46_23_c25;
   bh2587_w46_31_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_c25(0);
   bh2587_w47_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_c25(1);
   bh2587_w48_23_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2981: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2981_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_copy2982_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2981_Out0_copy2982_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2983_In0_c25 <= "" & bh2587_w47_22_c25 & bh2587_w47_20_c25 & bh2587_w47_18_c25 & bh2587_w47_16_c25 & bh2587_w47_15_c25 & bh2587_w47_17_c25;
   bh2587_w47_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_c25(0);
   bh2587_w48_24_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_c25(1);
   bh2587_w49_20_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2983: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2983_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_copy2984_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2983_Out0_copy2984_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid2985_In0_c25 <= "" & bh2587_w47_19_c25 & bh2587_w47_21_c25 & bh2587_w47_23_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid2985_In1_c25 <= "" & bh2587_w48_21_c25 & bh2587_w48_19_c25;
   bh2587_w47_28_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_c25(0);
   bh2587_w48_25_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_c25(1);
   bh2587_w49_21_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid2985: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid2985_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid2985_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_copy2986_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid2985_Out0_copy2986_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2987_In0_c25 <= "" & bh2587_w48_17_c25 & bh2587_w48_9_c25 & bh2587_w48_15_c25 & bh2587_w48_16_c25 & bh2587_w48_18_c25 & bh2587_w48_20_c25;
   bh2587_w48_26_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_c25(0);
   bh2587_w49_22_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_c25(1);
   bh2587_w50_18_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2987: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2987_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_copy2988_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2987_Out0_copy2988_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2989_In0_c25 <= "" & bh2587_w49_18_c25 & bh2587_w49_16_c25 & bh2587_w49_15_c25 & bh2587_w49_14_c25 & "0" & "0";
   bh2587_w49_23_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_c25(0);
   bh2587_w50_19_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_c25(1);
   bh2587_w51_15_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2989: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2989_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_copy2990_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2989_Out0_copy2990_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2991_In0_c25 <= "" & bh2587_w49_13_c25 & bh2587_w49_6_c25 & bh2587_w49_17_c25 & bh2587_w49_19_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2991_In1_c25 <= "" & bh2587_w50_17_c25;
   bh2587_w49_24_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_c25(0);
   bh2587_w50_20_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_c25(1);
   bh2587_w51_16_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2991: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2991_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2991_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_copy2992_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2991_Out0_copy2992_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2993_In0_c25 <= "" & bh2587_w50_11_c25 & bh2587_w50_12_c25 & bh2587_w50_13_c25 & bh2587_w50_14_c25 & bh2587_w50_15_c25 & bh2587_w50_16_c25;
   bh2587_w50_21_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_c25(0);
   bh2587_w51_17_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_c25(1);
   bh2587_w52_15_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2993: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2993_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_copy2994_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2993_Out0_copy2994_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2995_In0_c25 <= "" & bh2587_w51_9_c25 & bh2587_w51_10_c25 & bh2587_w51_11_c25 & bh2587_w51_12_c25 & bh2587_w51_13_c25 & bh2587_w51_14_c25;
   bh2587_w51_18_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_c25(0);
   bh2587_w52_16_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_c25(1);
   bh2587_w53_11_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2995: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2995_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_copy2996_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2995_Out0_copy2996_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid2997_In0_c25 <= "" & bh2587_w52_9_c25 & bh2587_w52_10_c25 & bh2587_w52_11_c25 & bh2587_w52_12_c25 & bh2587_w52_13_c25 & bh2587_w52_14_c25;
   bh2587_w52_17_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_c25(0);
   bh2587_w53_12_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_c25(1);
   bh2587_w54_10_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid2997: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid2997_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_copy2998_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid2997_Out0_copy2998_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In0_c25 <= "" & bh2587_w53_6_c25 & bh2587_w53_7_c25 & bh2587_w53_8_c25 & bh2587_w53_9_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In1_c24 <= "" & bh2587_w54_6_c24;
   bh2587_w53_13_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_c25(0);
   bh2587_w54_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_c25(1);
   bh2587_w55_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid2999: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid2999_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_copy3000_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid2999_Out0_copy3000_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3001_In0_c25 <= "" & bh2587_w54_7_c25 & bh2587_w54_8_c25 & bh2587_w54_9_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3001_In1_c25 <= "" & bh2587_w55_6_c25 & bh2587_w55_7_c25;
   bh2587_w54_12_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_c25(0);
   bh2587_w55_10_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_c25(1);
   bh2587_w56_8_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3001: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3001_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3001_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_copy3002_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3001_Out0_copy3002_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In0_c25 <= "" & bh2587_w56_4_c25 & bh2587_w56_5_c25 & bh2587_w56_6_c25 & bh2587_w56_7_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c0 <= "" & "0";
   bh2587_w56_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_c25(0);
   bh2587_w57_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_c25(1);
   bh2587_w58_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3003: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3003_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_copy3004_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3003_Out0_copy3004_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3005_In0_c25 <= "" & bh2587_w57_4_c25 & bh2587_w57_5_c25 & bh2587_w57_6_c25;
   bh2587_w57_8_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_c25(0);
   bh2587_w58_8_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3005: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3005_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_copy3006_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3005_Out0_copy3006_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3007_In0_c25 <= "" & bh2587_w58_4_c25 & bh2587_w58_5_c25 & bh2587_w58_6_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3007_In1_c25 <= "" & bh2587_w59_3_c25 & bh2587_w59_4_c25;
   bh2587_w58_9_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_c25(0);
   bh2587_w59_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_c25(1);
   bh2587_w60_6_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3007: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3007_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3007_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_copy3008_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3007_Out0_copy3008_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3009_In0_c25 <= "" & bh2587_w60_3_c25 & bh2587_w60_4_c25 & bh2587_w60_5_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3009_In1_c25 <= "" & bh2587_w61_2_c25 & bh2587_w61_3_c25;
   bh2587_w60_7_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_c25(0);
   bh2587_w61_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_c25(1);
   bh2587_w62_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3009: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3009_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3009_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_copy3010_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3009_Out0_copy3010_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3011_In0_c25 <= "" & bh2587_w62_3_c25 & bh2587_w62_4_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3011_In1_c25 <= "" & bh2587_w63_2_c25 & bh2587_w63_3_c25;
   bh2587_w62_6_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_c25(0);
   bh2587_w63_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_c25(1);
   bh2587_w64_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3011: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3011_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3011_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_copy3012_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3011_Out0_copy3012_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3013_In0_c25 <= "" & bh2587_w64_3_c25 & bh2587_w64_4_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3013_In1_c25 <= "" & bh2587_w65_2_c25 & bh2587_w65_3_c25;
   bh2587_w64_6_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_c25(0);
   bh2587_w65_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_c25(1);
   bh2587_w66_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3013: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3013_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3013_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_copy3014_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3013_Out0_copy3014_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3015_In0_c25 <= "" & bh2587_w66_3_c25 & bh2587_w66_4_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3015_In1_c25 <= "" & bh2587_w67_2_c25 & bh2587_w67_3_c25;
   bh2587_w66_6_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_c25(0);
   bh2587_w67_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_c25(1);
   bh2587_w68_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3015: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3015_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3015_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_copy3016_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3015_Out0_copy3016_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3017_In0_c25 <= "" & bh2587_w68_3_c25 & bh2587_w68_4_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3017_In1_c25 <= "" & bh2587_w69_2_c25 & bh2587_w69_3_c25;
   bh2587_w68_6_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_c25(0);
   bh2587_w69_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_c25(1);
   bh2587_w70_4_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3017: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3017_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3017_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_copy3018_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3017_Out0_copy3018_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3019_In0_c25 <= "" & bh2587_w70_2_c25 & bh2587_w70_3_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3019_In1_c25 <= "" & bh2587_w71_2_c25;
   bh2587_w70_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_c25(0);
   bh2587_w71_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_c25(1);
   bh2587_w72_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3019: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3019_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3019_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_copy3020_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3019_Out0_copy3020_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3021_In0_c25 <= "" & bh2587_w72_2_c25 & bh2587_w72_3_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3021_In1_c25 <= "" & bh2587_w73_2_c25;
   bh2587_w72_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_c25(0);
   bh2587_w73_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_c25(1);
   bh2587_w74_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3021: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3021_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3021_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_copy3022_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3021_Out0_copy3022_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3023_In0_c25 <= "" & bh2587_w74_2_c25 & bh2587_w74_3_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3023_In1_c25 <= "" & bh2587_w75_2_c25;
   bh2587_w74_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_c25(0);
   bh2587_w75_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_c25(1);
   bh2587_w76_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3023: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3023_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3023_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_copy3024_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3023_Out0_copy3024_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3025_In0_c25 <= "" & bh2587_w76_0_c25 & bh2587_w76_1_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3025_In1_c25 <= "" & bh2587_w77_0_c25;
   bh2587_w76_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_c25(0);
   bh2587_w77_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_c25(1);
   bh2587_w78_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3025: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3025_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3025_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_copy3026_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3025_Out0_copy3026_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3027_In0_c25 <= "" & bh2587_w38_4_c25 & "0" & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3027_In1_c25 <= "" & bh2587_w39_34_c25 & bh2587_w39_35_c25;
   bh2587_w38_5_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_c25(0);
   bh2587_w39_36_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_c25(1);
   bh2587_w40_30_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3027: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3027_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3027_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_copy3028_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3027_Out0_copy3028_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3029_In0_c25 <= "" & bh2587_w40_27_c25 & bh2587_w40_28_c25 & bh2587_w40_29_c25;
   bh2587_w40_31_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_c25(0);
   bh2587_w41_34_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3029: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3029_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_copy3030_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3029_Out0_copy3030_c25; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid3032_bh2587_uid3033_In0_c25 <= "" & bh2587_w41_29_c25 & bh2587_w41_30_c25 & bh2587_w41_31_c25 & bh2587_w41_32_c25 & bh2587_w41_33_c25;
   bh2587_w41_35_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_c25(0);
   bh2587_w42_38_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_c25(1);
   bh2587_w43_38_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_c25(2);
   Compressor_5_3_Freq300_uid3032_uid3033: Compressor_5_3_Freq300_uid3032
      port map ( X0 => Compressor_5_3_Freq300_uid3032_bh2587_uid3033_In0_c25,
                 R => Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_copy3034_c25);
   Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3033_Out0_copy3034_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid3035_In0_c25 <= "" & bh2587_w42_32_c25 & bh2587_w42_33_c25 & bh2587_w42_34_c25 & bh2587_w42_35_c25 & bh2587_w42_36_c25 & bh2587_w42_37_c25;
   bh2587_w42_39_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_c25(0);
   bh2587_w43_39_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_c25(1);
   bh2587_w44_36_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid3035: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid3035_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_copy3036_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3035_Out0_copy3036_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid3037_In0_c25 <= "" & bh2587_w43_31_c25 & bh2587_w43_32_c25 & bh2587_w43_33_c25 & bh2587_w43_34_c25 & bh2587_w43_35_c25 & bh2587_w43_36_c25;
   bh2587_w43_40_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_c25(0);
   bh2587_w44_37_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_c25(1);
   bh2587_w45_34_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid3037: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid3037_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_copy3038_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3037_Out0_copy3038_c25; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid3032_bh2587_uid3039_In0_c25 <= "" & bh2587_w44_31_c25 & bh2587_w44_32_c25 & bh2587_w44_33_c25 & bh2587_w44_34_c25 & bh2587_w44_35_c25;
   bh2587_w44_38_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_c25(0);
   bh2587_w45_35_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_c25(1);
   bh2587_w46_32_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_c25(2);
   Compressor_5_3_Freq300_uid3032_uid3039: Compressor_5_3_Freq300_uid3032
      port map ( X0 => Compressor_5_3_Freq300_uid3032_bh2587_uid3039_In0_c25,
                 R => Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_copy3040_c25);
   Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_c25 <= Compressor_5_3_Freq300_uid3032_bh2587_uid3039_Out0_copy3040_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid3041_In0_c25 <= "" & bh2587_w45_28_c25 & bh2587_w45_29_c25 & bh2587_w45_30_c25 & bh2587_w45_31_c25 & bh2587_w45_32_c25 & bh2587_w45_33_c25;
   bh2587_w45_36_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_c25(0);
   bh2587_w46_33_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_c25(1);
   bh2587_w47_29_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid3041: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid3041_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_copy3042_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3041_Out0_copy3042_c25; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid2838_bh2587_uid3043_In0_c25 <= "" & bh2587_w46_25_c25 & bh2587_w46_27_c25 & bh2587_w46_28_c25 & bh2587_w46_29_c25 & bh2587_w46_30_c25 & bh2587_w46_31_c25;
   bh2587_w46_34_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_c25(0);
   bh2587_w47_30_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_c25(1);
   bh2587_w48_27_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_c25(2);
   Compressor_6_3_Freq300_uid2838_uid3043: Compressor_6_3_Freq300_uid2838
      port map ( X0 => Compressor_6_3_Freq300_uid2838_bh2587_uid3043_In0_c25,
                 R => Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_copy3044_c25);
   Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_c25 <= Compressor_6_3_Freq300_uid2838_bh2587_uid3043_Out0_copy3044_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3045_In0_c25 <= "" & bh2587_w47_24_c25 & bh2587_w47_25_c25 & bh2587_w47_26_c25 & bh2587_w47_27_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3045_In1_c25 <= "" & bh2587_w48_22_c25;
   bh2587_w47_31_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_c25(0);
   bh2587_w48_28_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_c25(1);
   bh2587_w49_25_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3045: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3045_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3045_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_copy3046_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3045_Out0_copy3046_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3047_In0_c25 <= "" & bh2587_w48_23_c25 & bh2587_w48_24_c25 & bh2587_w48_25_c25 & bh2587_w48_26_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3047_In1_c25 <= "" & bh2587_w49_20_c25;
   bh2587_w48_29_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_c25(0);
   bh2587_w49_26_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_c25(1);
   bh2587_w50_22_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3047: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3047_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3047_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_copy3048_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3047_Out0_copy3048_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3049_In0_c25 <= "" & bh2587_w49_21_c25 & bh2587_w49_22_c25 & bh2587_w49_23_c25 & bh2587_w49_24_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3049_In1_c25 <= "" & bh2587_w50_18_c25;
   bh2587_w49_27_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_c25(0);
   bh2587_w50_23_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_c25(1);
   bh2587_w51_19_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3049: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3049_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3049_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_copy3050_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3049_Out0_copy3050_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3051_In0_c25 <= "" & bh2587_w50_19_c25 & bh2587_w50_20_c25 & bh2587_w50_21_c25;
   bh2587_w50_24_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_c25(0);
   bh2587_w51_20_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3051: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3051_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_copy3052_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3051_Out0_copy3052_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In0_c25 <= "" & bh2587_w51_15_c25 & bh2587_w51_16_c25 & bh2587_w51_17_c25 & bh2587_w51_18_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c0 <= "" & "0";
   bh2587_w51_21_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_c25(0);
   bh2587_w52_18_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_c25(1);
   bh2587_w53_14_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3053: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3053_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_copy3054_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3053_Out0_copy3054_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3055_In0_c25 <= "" & bh2587_w52_15_c25 & bh2587_w52_16_c25 & bh2587_w52_17_c25;
   bh2587_w52_19_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_c25(0);
   bh2587_w53_15_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3055: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3055_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_copy3056_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3055_Out0_copy3056_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In0_c25 <= "" & bh2587_w53_10_c25 & bh2587_w53_11_c25 & bh2587_w53_12_c25 & bh2587_w53_13_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c0 <= "" & "0";
   bh2587_w53_16_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_c25(0);
   bh2587_w54_13_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_c25(1);
   bh2587_w55_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3057: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3057_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_copy3058_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3057_Out0_copy3058_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3059_In0_c25 <= "" & bh2587_w54_10_c25 & bh2587_w54_11_c25 & bh2587_w54_12_c25;
   bh2587_w54_14_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_c25(0);
   bh2587_w55_12_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3059: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3059_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_copy3060_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3059_Out0_copy3060_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3061_In0_c25 <= "" & bh2587_w55_8_c25 & bh2587_w55_9_c25 & bh2587_w55_10_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3061_In1_c25 <= "" & bh2587_w56_8_c25 & bh2587_w56_9_c25;
   bh2587_w55_13_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_c25(0);
   bh2587_w56_10_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_c25(1);
   bh2587_w57_9_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3061: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3061_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3061_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_copy3062_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3061_Out0_copy3062_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3063_In0_c25 <= "" & bh2587_w57_7_c25 & bh2587_w57_8_c25 & "0";
   bh2587_w57_10_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_c25(0);
   bh2587_w58_10_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3063: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3063_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_copy3064_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3063_Out0_copy3064_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3065_In0_c25 <= "" & bh2587_w58_7_c25 & bh2587_w58_8_c25 & bh2587_w58_9_c25;
   bh2587_w58_11_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_c25(0);
   bh2587_w59_6_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3065: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3065_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_copy3066_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3065_Out0_copy3066_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3067_In0_c25 <= "" & bh2587_w60_6_c25 & bh2587_w60_7_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3067_In1_c25 <= "" & bh2587_w61_4_c25;
   bh2587_w60_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_c25(0);
   bh2587_w61_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_c25(1);
   bh2587_w62_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3067: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3067_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3067_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_copy3068_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3067_Out0_copy3068_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3069_In0_c25 <= "" & bh2587_w62_5_c25 & bh2587_w62_6_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3069_In1_c25 <= "" & bh2587_w63_4_c25;
   bh2587_w62_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_c25(0);
   bh2587_w63_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_c25(1);
   bh2587_w64_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3069: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3069_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3069_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_copy3070_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3069_Out0_copy3070_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3071_In0_c25 <= "" & bh2587_w64_5_c25 & bh2587_w64_6_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3071_In1_c25 <= "" & bh2587_w65_4_c25;
   bh2587_w64_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_c25(0);
   bh2587_w65_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_c25(1);
   bh2587_w66_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3071: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3071_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3071_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_copy3072_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3071_Out0_copy3072_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3073_In0_c25 <= "" & bh2587_w66_5_c25 & bh2587_w66_6_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3073_In1_c25 <= "" & bh2587_w67_4_c25;
   bh2587_w66_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_c25(0);
   bh2587_w67_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_c25(1);
   bh2587_w68_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3073: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3073_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3073_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_copy3074_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3073_Out0_copy3074_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3075_In0_c25 <= "" & bh2587_w68_5_c25 & bh2587_w68_6_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3075_In1_c25 <= "" & bh2587_w69_4_c25;
   bh2587_w68_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_c25(0);
   bh2587_w69_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_c25(1);
   bh2587_w70_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3075: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3075_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3075_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_copy3076_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3075_Out0_copy3076_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3077_In0_c25 <= "" & bh2587_w70_4_c25 & bh2587_w70_5_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3077_In1_c25 <= "" & bh2587_w71_3_c25;
   bh2587_w70_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_c25(0);
   bh2587_w71_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_c25(1);
   bh2587_w72_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3077: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3077_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3077_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_copy3078_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3077_Out0_copy3078_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3079_In0_c25 <= "" & bh2587_w72_4_c25 & bh2587_w72_5_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3079_In1_c25 <= "" & bh2587_w73_3_c25;
   bh2587_w72_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_c25(0);
   bh2587_w73_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_c25(1);
   bh2587_w74_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3079: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3079_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3079_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_copy3080_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3079_Out0_copy3080_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3081_In0_c25 <= "" & bh2587_w74_4_c25 & bh2587_w74_5_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3081_In1_c25 <= "" & bh2587_w75_3_c25;
   bh2587_w74_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_c25(0);
   bh2587_w75_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_c25(1);
   bh2587_w76_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3081: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3081_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3081_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_copy3082_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3081_Out0_copy3082_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3083_In0_c25 <= "" & bh2587_w76_2_c25 & bh2587_w76_3_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3083_In1_c25 <= "" & bh2587_w77_1_c25;
   bh2587_w76_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_c25(0);
   bh2587_w77_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_c25(1);
   bh2587_w78_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3083: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3083_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3083_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_copy3084_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3083_Out0_copy3084_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3085_In0_c25 <= "" & bh2587_w78_0_c25 & bh2587_w78_1_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3085_In1_c25 <= "" & bh2587_w79_0_c25;
   bh2587_w78_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_c25(0);
   bh2587_w79_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_c25(1);
   bh2587_w80_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3085: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3085_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3085_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_copy3086_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3085_Out0_copy3086_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3087_In0_c25 <= "" & bh2587_w40_30_c25 & bh2587_w40_31_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3087_In1_c25 <= "" & bh2587_w41_34_c25 & bh2587_w41_35_c25;
   bh2587_w40_32_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_c25(0);
   bh2587_w41_36_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_c25(1);
   bh2587_w42_40_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3087: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3087_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3087_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_copy3088_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3087_Out0_copy3088_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3089_In0_c25 <= "" & bh2587_w42_38_c25 & bh2587_w42_39_c25 & "0";
   bh2587_w42_41_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_c25(0);
   bh2587_w43_41_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3089: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3089_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_copy3090_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3089_Out0_copy3090_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In0_c25 <= "" & bh2587_w43_37_c25 & bh2587_w43_38_c25 & bh2587_w43_39_c25 & bh2587_w43_40_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c0 <= "" & "0";
   bh2587_w43_42_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_c25(0);
   bh2587_w44_39_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_c25(1);
   bh2587_w45_37_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3091: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3091_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_copy3092_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3091_Out0_copy3092_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3093_In0_c25 <= "" & bh2587_w44_36_c25 & bh2587_w44_37_c25 & bh2587_w44_38_c25;
   bh2587_w44_40_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_c25(0);
   bh2587_w45_38_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3093: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3093_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_copy3094_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3093_Out0_copy3094_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3095_In0_c25 <= "" & bh2587_w45_34_c25 & bh2587_w45_35_c25 & bh2587_w45_36_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3095_In1_c25 <= "" & bh2587_w46_32_c25 & bh2587_w46_33_c25;
   bh2587_w45_39_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_c25(0);
   bh2587_w46_35_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_c25(1);
   bh2587_w47_32_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3095: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3095_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3095_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_copy3096_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3095_Out0_copy3096_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In0_c25 <= "" & bh2587_w47_28_c25 & bh2587_w47_29_c25 & bh2587_w47_30_c25 & bh2587_w47_31_c25;
   Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c0 <= "" & "0";
   bh2587_w47_33_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_c25(0);
   bh2587_w48_30_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_c25(1);
   bh2587_w49_28_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3097: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3097_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_copy3098_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3097_Out0_copy3098_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3099_In0_c25 <= "" & bh2587_w48_27_c25 & bh2587_w48_28_c25 & bh2587_w48_29_c25;
   bh2587_w48_31_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_c25(0);
   bh2587_w49_29_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3099: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3099_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_copy3100_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3099_Out0_copy3100_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3101_In0_c25 <= "" & bh2587_w49_25_c25 & bh2587_w49_26_c25 & bh2587_w49_27_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3101_In1_c25 <= "" & bh2587_w50_22_c25 & bh2587_w50_23_c25;
   bh2587_w49_30_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_c25(0);
   bh2587_w50_25_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_c25(1);
   bh2587_w51_22_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3101: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3101_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3101_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_copy3102_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3101_Out0_copy3102_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3103_In0_c25 <= "" & bh2587_w51_19_c25 & bh2587_w51_20_c25 & bh2587_w51_21_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3103_In1_c25 <= "" & bh2587_w52_18_c25 & bh2587_w52_19_c25;
   bh2587_w51_23_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_c25(0);
   bh2587_w52_20_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_c25(1);
   bh2587_w53_17_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3103: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3103_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3103_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_copy3104_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3103_Out0_copy3104_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3105_In0_c25 <= "" & bh2587_w53_14_c25 & bh2587_w53_15_c25 & bh2587_w53_16_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3105_In1_c25 <= "" & bh2587_w54_13_c25 & bh2587_w54_14_c25;
   bh2587_w53_18_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_c25(0);
   bh2587_w54_15_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_c25(1);
   bh2587_w55_14_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3105: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3105_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3105_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_copy3106_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3105_Out0_copy3106_c25; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3107_In0_c25 <= "" & bh2587_w55_11_c25 & bh2587_w55_12_c25 & bh2587_w55_13_c25;
   bh2587_w55_15_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_c25(0);
   bh2587_w56_11_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_c25(1);
   Compressor_3_2_Freq300_uid2834_uid3107: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3107_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_copy3108_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_c25 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3107_Out0_copy3108_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3109_In0_c25 <= "" & bh2587_w57_9_c25 & bh2587_w57_10_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3109_In1_c25 <= "" & bh2587_w58_10_c25 & bh2587_w58_11_c25;
   bh2587_w57_11_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_c25(0);
   bh2587_w58_12_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_c25(1);
   bh2587_w59_7_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_c25(2);
   Compressor_23_3_Freq300_uid2830_uid3109: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3109_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3109_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_copy3110_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_c25 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3109_Out0_copy3110_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3111_In0_c25 <= "" & bh2587_w59_5_c25 & bh2587_w59_6_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3111_In1_c25 <= "" & bh2587_w60_8_c25;
   bh2587_w59_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_c25(0);
   bh2587_w60_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_c25(1);
   bh2587_w61_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3111: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3111_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3111_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_copy3112_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3111_Out0_copy3112_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3113_In0_c25 <= "" & bh2587_w62_7_c25 & bh2587_w62_8_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3113_In1_c25 <= "" & bh2587_w63_5_c25;
   bh2587_w62_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_c25(0);
   bh2587_w63_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_c25(1);
   bh2587_w64_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3113: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3113_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3113_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_copy3114_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3113_Out0_copy3114_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3115_In0_c25 <= "" & bh2587_w64_7_c25 & bh2587_w64_8_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3115_In1_c25 <= "" & bh2587_w65_5_c25;
   bh2587_w64_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_c25(0);
   bh2587_w65_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_c25(1);
   bh2587_w66_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3115: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3115_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3115_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_copy3116_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3115_Out0_copy3116_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3117_In0_c25 <= "" & bh2587_w66_7_c25 & bh2587_w66_8_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3117_In1_c25 <= "" & bh2587_w67_5_c25;
   bh2587_w66_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_c25(0);
   bh2587_w67_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_c25(1);
   bh2587_w68_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3117: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3117_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3117_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_copy3118_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3117_Out0_copy3118_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3119_In0_c25 <= "" & bh2587_w68_7_c25 & bh2587_w68_8_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3119_In1_c25 <= "" & bh2587_w69_5_c25;
   bh2587_w68_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_c25(0);
   bh2587_w69_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_c25(1);
   bh2587_w70_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3119: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3119_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3119_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_copy3120_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3119_Out0_copy3120_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3121_In0_c25 <= "" & bh2587_w70_6_c25 & bh2587_w70_7_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3121_In1_c25 <= "" & bh2587_w71_4_c25;
   bh2587_w70_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_c25(0);
   bh2587_w71_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_c25(1);
   bh2587_w72_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3121: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3121_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3121_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_copy3122_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3121_Out0_copy3122_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3123_In0_c25 <= "" & bh2587_w72_6_c25 & bh2587_w72_7_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3123_In1_c25 <= "" & bh2587_w73_4_c25;
   bh2587_w72_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_c25(0);
   bh2587_w73_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_c25(1);
   bh2587_w74_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3123: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3123_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3123_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_copy3124_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3123_Out0_copy3124_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3125_In0_c25 <= "" & bh2587_w74_6_c25 & bh2587_w74_7_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3125_In1_c25 <= "" & bh2587_w75_4_c25;
   bh2587_w74_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_c25(0);
   bh2587_w75_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_c25(1);
   bh2587_w76_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3125: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3125_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3125_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_copy3126_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3125_Out0_copy3126_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3127_In0_c25 <= "" & bh2587_w76_4_c25 & bh2587_w76_5_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3127_In1_c25 <= "" & bh2587_w77_2_c25;
   bh2587_w76_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_c25(0);
   bh2587_w77_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_c25(1);
   bh2587_w78_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3127: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3127_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3127_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_copy3128_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3127_Out0_copy3128_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3129_In0_c25 <= "" & bh2587_w78_2_c25 & bh2587_w78_3_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3129_In1_c25 <= "" & bh2587_w79_1_c25;
   bh2587_w78_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_c25(0);
   bh2587_w79_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_c25(1);
   bh2587_w80_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3129: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3129_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3129_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_copy3130_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3129_Out0_copy3130_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3131_In0_c25 <= "" & bh2587_w80_0_c25 & bh2587_w80_1_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3131_In1_c25 <= "" & bh2587_w81_0_c25;
   bh2587_w80_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_c25(0);
   bh2587_w81_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_c25(1);
   bh2587_w82_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3131: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3131_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3131_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_copy3132_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3131_Out0_copy3132_c25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3133_In0_c25 <= "" & bh2587_w42_40_c25 & bh2587_w42_41_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3133_In1_c25 <= "" & bh2587_w43_41_c25 & bh2587_w43_42_c25;
   bh2587_w42_42_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_c26(0);
   bh2587_w43_43_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_c26(1);
   bh2587_w44_41_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_c26(2);
   Compressor_23_3_Freq300_uid2830_uid3133: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3133_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3133_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_copy3134_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3133_Out0_copy3134_c26; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid2834_bh2587_uid3135_In0_c25 <= "" & bh2587_w44_39_c25 & bh2587_w44_40_c25 & "0";
   bh2587_w44_42_c26 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_c26(0);
   bh2587_w45_40_c26 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_c26(1);
   Compressor_3_2_Freq300_uid2834_uid3135: Compressor_3_2_Freq300_uid2834
      port map ( X0 => Compressor_3_2_Freq300_uid2834_bh2587_uid3135_In0_c25,
                 R => Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_copy3136_c25);
   Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_c26 <= Compressor_3_2_Freq300_uid2834_bh2587_uid3135_Out0_copy3136_c26; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3137_In0_c25 <= "" & bh2587_w45_37_c25 & bh2587_w45_38_c25 & bh2587_w45_39_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3137_In1_c25 <= "" & bh2587_w46_34_c25 & bh2587_w46_35_c25;
   bh2587_w45_41_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_c26(0);
   bh2587_w46_36_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_c26(1);
   bh2587_w47_34_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_c26(2);
   Compressor_23_3_Freq300_uid2830_uid3137: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3137_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3137_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_copy3138_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3137_Out0_copy3138_c26; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3139_In0_c25 <= "" & bh2587_w47_32_c25 & bh2587_w47_33_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3139_In1_c25 <= "" & bh2587_w48_30_c25 & bh2587_w48_31_c25;
   bh2587_w47_35_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_c26(0);
   bh2587_w48_32_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_c26(1);
   bh2587_w49_31_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_c26(2);
   Compressor_23_3_Freq300_uid2830_uid3139: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3139_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3139_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_copy3140_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3139_Out0_copy3140_c26; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3141_In0_c25 <= "" & bh2587_w49_28_c25 & bh2587_w49_29_c25 & bh2587_w49_30_c25;
   Compressor_23_3_Freq300_uid2830_bh2587_uid3141_In1_c25 <= "" & bh2587_w50_24_c25 & bh2587_w50_25_c25;
   bh2587_w49_32_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_c26(0);
   bh2587_w50_26_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_c26(1);
   bh2587_w51_24_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_c26(2);
   Compressor_23_3_Freq300_uid2830_uid3141: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3141_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3141_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_copy3142_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3141_Out0_copy3142_c26; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3143_In0_c25 <= "" & bh2587_w51_22_c25 & bh2587_w51_23_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3143_In1_c25 <= "" & bh2587_w52_20_c25;
   bh2587_w51_25_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_c26(0);
   bh2587_w52_21_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_c26(1);
   bh2587_w53_19_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_c26(2);
   Compressor_14_3_Freq300_uid2848_uid3143: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3143_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3143_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_copy3144_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3143_Out0_copy3144_c26; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3145_In0_c25 <= "" & bh2587_w53_17_c25 & bh2587_w53_18_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3145_In1_c25 <= "" & bh2587_w54_15_c25;
   bh2587_w53_20_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_c26(0);
   bh2587_w54_16_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_c26(1);
   bh2587_w55_16_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_c26(2);
   Compressor_14_3_Freq300_uid2848_uid3145: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3145_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3145_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_copy3146_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_c26 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3145_Out0_copy3146_c26; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid2830_bh2587_uid3147_In0_c25 <= "" & bh2587_w55_14_c25 & bh2587_w55_15_c25 & "0";
   Compressor_23_3_Freq300_uid2830_bh2587_uid3147_In1_c25 <= "" & bh2587_w56_10_c25 & bh2587_w56_11_c25;
   bh2587_w55_17_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_c26(0);
   bh2587_w56_12_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_c26(1);
   bh2587_w57_12_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_c26(2);
   Compressor_23_3_Freq300_uid2830_uid3147: Compressor_23_3_Freq300_uid2830
      port map ( X0 => Compressor_23_3_Freq300_uid2830_bh2587_uid3147_In0_c25,
                 X1 => Compressor_23_3_Freq300_uid2830_bh2587_uid3147_In1_c25,
                 R => Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_copy3148_c25);
   Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_c26 <= Compressor_23_3_Freq300_uid2830_bh2587_uid3147_Out0_copy3148_c26; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3149_In0_c25 <= "" & bh2587_w59_7_c25 & bh2587_w59_8_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3149_In1_c25 <= "" & bh2587_w60_9_c25;
   bh2587_w59_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_c25(0);
   bh2587_w60_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_c25(1);
   bh2587_w61_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3149: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3149_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3149_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_copy3150_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3149_Out0_copy3150_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3151_In0_c25 <= "" & bh2587_w61_5_c25 & bh2587_w61_6_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3151_In1_c25 <= "" & bh2587_w62_9_c25;
   bh2587_w61_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_c25(0);
   bh2587_w62_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_c25(1);
   bh2587_w63_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3151: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3151_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3151_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_copy3152_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3151_Out0_copy3152_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3153_In0_c25 <= "" & bh2587_w64_9_c25 & bh2587_w64_10_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3153_In1_c25 <= "" & bh2587_w65_6_c25;
   bh2587_w64_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_c25(0);
   bh2587_w65_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_c25(1);
   bh2587_w66_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3153: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3153_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3153_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_copy3154_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3153_Out0_copy3154_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3155_In0_c25 <= "" & bh2587_w66_9_c25 & bh2587_w66_10_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3155_In1_c25 <= "" & bh2587_w67_6_c25;
   bh2587_w66_12_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_c25(0);
   bh2587_w67_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_c25(1);
   bh2587_w68_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3155: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3155_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3155_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_copy3156_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3155_Out0_copy3156_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3157_In0_c25 <= "" & bh2587_w68_9_c25 & bh2587_w68_10_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3157_In1_c25 <= "" & bh2587_w69_6_c25;
   bh2587_w68_12_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_c25(0);
   bh2587_w69_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_c25(1);
   bh2587_w70_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3157: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3157_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3157_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_copy3158_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3157_Out0_copy3158_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3159_In0_c25 <= "" & bh2587_w70_8_c25 & bh2587_w70_9_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3159_In1_c25 <= "" & bh2587_w71_5_c25;
   bh2587_w70_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_c25(0);
   bh2587_w71_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_c25(1);
   bh2587_w72_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3159: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3159_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3159_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_copy3160_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3159_Out0_copy3160_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3161_In0_c25 <= "" & bh2587_w72_8_c25 & bh2587_w72_9_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3161_In1_c25 <= "" & bh2587_w73_5_c25;
   bh2587_w72_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_c25(0);
   bh2587_w73_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_c25(1);
   bh2587_w74_10_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3161: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3161_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3161_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_copy3162_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3161_Out0_copy3162_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3163_In0_c25 <= "" & bh2587_w74_8_c25 & bh2587_w74_9_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3163_In1_c25 <= "" & bh2587_w75_5_c25;
   bh2587_w74_11_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_c25(0);
   bh2587_w75_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_c25(1);
   bh2587_w76_8_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3163: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3163_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3163_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_copy3164_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3163_Out0_copy3164_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3165_In0_c25 <= "" & bh2587_w76_6_c25 & bh2587_w76_7_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3165_In1_c25 <= "" & bh2587_w77_3_c25;
   bh2587_w76_9_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_c25(0);
   bh2587_w77_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_c25(1);
   bh2587_w78_6_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3165: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3165_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3165_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_copy3166_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3165_Out0_copy3166_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3167_In0_c25 <= "" & bh2587_w78_4_c25 & bh2587_w78_5_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3167_In1_c25 <= "" & bh2587_w79_2_c25;
   bh2587_w78_7_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_c25(0);
   bh2587_w79_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_c25(1);
   bh2587_w80_4_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3167: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3167_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3167_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_copy3168_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3167_Out0_copy3168_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3169_In0_c25 <= "" & bh2587_w80_2_c25 & bh2587_w80_3_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3169_In1_c25 <= "" & bh2587_w81_1_c25;
   bh2587_w80_5_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_c25(0);
   bh2587_w81_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_c25(1);
   bh2587_w82_2_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3169: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3169_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3169_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_copy3170_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3169_Out0_copy3170_c25; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid2848_bh2587_uid3171_In0_c25 <= "" & bh2587_w82_0_c25 & bh2587_w82_1_c25 & "0" & "0";
   Compressor_14_3_Freq300_uid2848_bh2587_uid3171_In1_c25 <= "" & bh2587_w83_0_c25;
   bh2587_w82_3_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_c25(0);
   bh2587_w83_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_c25(1);
   bh2587_w84_1_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_c25(2);
   Compressor_14_3_Freq300_uid2848_uid3171: Compressor_14_3_Freq300_uid2848
      port map ( X0 => Compressor_14_3_Freq300_uid2848_bh2587_uid3171_In0_c25,
                 X1 => Compressor_14_3_Freq300_uid2848_bh2587_uid3171_In1_c25,
                 R => Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_copy3172_c25);
   Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_c25 <= Compressor_14_3_Freq300_uid2848_bh2587_uid3171_Out0_copy3172_c25; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh2587_43_c26 <= bh2587_w43_43_c26 & bh2587_w42_42_c26 & bh2587_w41_36_c26 & bh2587_w40_32_c26 & bh2587_w39_36_c26 & bh2587_w38_5_c26 & bh2587_w37_3_c26 & bh2587_w36_2_c26 & bh2587_w35_0_c26 & bh2587_w34_0_c26 & bh2587_w33_0_c26 & bh2587_w32_0_c26 & bh2587_w31_0_c26 & bh2587_w30_0_c26 & bh2587_w29_0_c26 & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0";

   bitheapFinalAdd_bh2587_In0_c26 <= "0" & bh2587_w92_0_c26 & bh2587_w91_0_c26 & bh2587_w90_0_c26 & bh2587_w89_0_c26 & bh2587_w88_0_c26 & bh2587_w87_0_c26 & bh2587_w86_0_c26 & bh2587_w85_0_c26 & bh2587_w84_0_c26 & bh2587_w83_1_c26 & bh2587_w82_2_c26 & bh2587_w81_2_c26 & bh2587_w80_4_c26 & bh2587_w79_3_c26 & bh2587_w78_6_c26 & bh2587_w77_4_c26 & bh2587_w76_8_c26 & bh2587_w75_6_c26 & bh2587_w74_10_c26 & bh2587_w73_6_c26 & bh2587_w72_10_c26 & bh2587_w71_6_c26 & bh2587_w70_10_c26 & bh2587_w69_7_c26 & bh2587_w68_11_c26 & bh2587_w67_7_c26 & bh2587_w66_11_c26 & bh2587_w65_7_c26 & bh2587_w64_11_c26 & bh2587_w63_6_c26 & bh2587_w62_10_c26 & bh2587_w61_7_c26 & bh2587_w60_10_c26 & bh2587_w59_9_c26 & bh2587_w58_12_c26 & bh2587_w57_11_c26 & bh2587_w56_12_c26 & bh2587_w55_16_c26 & bh2587_w54_16_c26 & bh2587_w53_19_c26 & bh2587_w52_21_c26 & bh2587_w51_24_c26 & bh2587_w50_26_c26 & bh2587_w49_31_c26 & bh2587_w48_32_c26 & bh2587_w47_34_c26 & bh2587_w46_36_c26 & bh2587_w45_40_c26 & bh2587_w44_41_c26;
   bitheapFinalAdd_bh2587_In1_c26 <= "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & bh2587_w84_1_c26 & "0" & bh2587_w82_3_c26 & "0" & bh2587_w80_5_c26 & "0" & bh2587_w78_7_c26 & "0" & bh2587_w76_9_c26 & "0" & bh2587_w74_11_c26 & "0" & bh2587_w72_11_c26 & "0" & bh2587_w70_11_c26 & "0" & bh2587_w68_12_c26 & "0" & bh2587_w66_12_c26 & "0" & "0" & bh2587_w63_7_c26 & "0" & bh2587_w61_8_c26 & "0" & "0" & "0" & bh2587_w57_12_c26 & "0" & bh2587_w55_17_c26 & "0" & bh2587_w53_20_c26 & "0" & bh2587_w51_25_c26 & "0" & bh2587_w49_32_c26 & "0" & bh2587_w47_35_c26 & "0" & bh2587_w45_41_c26 & bh2587_w44_42_c26;
   bitheapFinalAdd_bh2587_Cin_c0 <= '0';

   bitheapFinalAdd_bh2587: IntAdder_50_Freq300_uid3174
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 Cin => bitheapFinalAdd_bh2587_Cin_c0,
                 X => bitheapFinalAdd_bh2587_In0_c26,
                 Y => bitheapFinalAdd_bh2587_In1_c26,
                 R => bitheapFinalAdd_bh2587_Out_c26);
   bitheapResult_bh2587_c26 <= bitheapFinalAdd_bh2587_Out_c26(48 downto 0) & tmp_bitheapResult_bh2587_43_c26;
   R <= bitheapResult_bh2587_c26(92 downto 45);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_57_Freq300_uid3177
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_57_Freq300_uid3177 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27 : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Y : in  std_logic_vector(56 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of IntAdder_57_Freq300_uid3177 is
signal Rtmp_c27 :  std_logic_vector(56 downto 0);
signal X_c21, X_c22, X_c23, X_c24, X_c25, X_c26, X_c27 :  std_logic_vector(56 downto 0);
signal Y_c27 :  std_logic_vector(56 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19, Cin_c20, Cin_c21, Cin_c22, Cin_c23, Cin_c24, Cin_c25, Cin_c26, Cin_c27 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               Cin_c19 <= Cin_c18;
            end if;
            if ce_20 = '1' then
               Cin_c20 <= Cin_c19;
            end if;
            if ce_21 = '1' then
               X_c21 <= X;
               Cin_c21 <= Cin_c20;
            end if;
            if ce_22 = '1' then
               X_c22 <= X_c21;
               Cin_c22 <= Cin_c21;
            end if;
            if ce_23 = '1' then
               X_c23 <= X_c22;
               Cin_c23 <= Cin_c22;
            end if;
            if ce_24 = '1' then
               X_c24 <= X_c23;
               Cin_c24 <= Cin_c23;
            end if;
            if ce_25 = '1' then
               X_c25 <= X_c24;
               Cin_c25 <= Cin_c24;
            end if;
            if ce_26 = '1' then
               X_c26 <= X_c25;
               Cin_c26 <= Cin_c25;
            end if;
            if ce_27 = '1' then
               X_c27 <= X_c26;
               Y_c27 <= Y;
               Cin_c27 <= Cin_c26;
            end if;
         end if;
      end process;
   Rtmp_c27 <= X_c27 + Y_c27 + Cin_c27;
   R <= Rtmp_c27;
end architecture;

--------------------------------------------------------------------------------
--                         Exp_11_52_Freq300_uid1481
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: ufixX_i XSign
-- Output signals: expY K

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Exp_11_52_Freq300_uid1481 is
    port (clk, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27 : in std_logic;
          ufixX_i : in  std_logic_vector(65 downto 0);
          XSign : in  std_logic;
          expY : out  std_logic_vector(56 downto 0);
          K : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of Exp_11_52_Freq300_uid1481 is
   component FixRealKCM_Freq300_uid1483 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(10 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid1510 is
      port ( clk, ce_18 : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             R : out  std_logic_vector(66 downto 0)   );
   end component;

   component IntAdder_56_Freq300_uid1523 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19 : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component FixFunctionByTable_Freq300_uid1525 is
      port ( clk, ce_20 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(56 downto 0)   );
   end component;

   component FixFunctionByPiecewisePoly_Freq300_uid1534 is
      port ( clk, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             X : in  std_logic_vector(35 downto 0);
             Y : out  std_logic_vector(35 downto 0)   );
   end component;

   component IntAdder_47_Freq300_uid2583 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24 : in std_logic;
             X : in  std_logic_vector(46 downto 0);
             Y : in  std_logic_vector(46 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(46 downto 0)   );
   end component;

   component IntMultiplier_46x47_48_Freq300_uid2585 is
      port ( clk, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
             X : in  std_logic_vector(45 downto 0);
             Y : in  std_logic_vector(46 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_57_Freq300_uid3177 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27 : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Y : in  std_logic_vector(56 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(56 downto 0)   );
   end component;

signal ufixX_c17 :  unsigned(9+56 downto 0);
signal xMulIn_c17 :  unsigned(9+3 downto 0);
signal absK_c17, absK_c18 :  std_logic_vector(10 downto 0);
signal minusAbsK_c18 :  std_logic_vector(11 downto 0);
signal absKLog2_c18 :  std_logic_vector(66 downto 0);
signal subOp1_c17 :  std_logic_vector(55 downto 0);
signal subOp2_c18 :  std_logic_vector(55 downto 0);
signal Y_c19 :  std_logic_vector(55 downto 0);
signal A_c19 :  std_logic_vector(9 downto 0);
signal Z_c19 :  std_logic_vector(45 downto 0);
signal expA_c20 :  std_logic_vector(56 downto 0);
signal Ztrunc_c19 :  std_logic_vector(35 downto 0);
signal expZmZm1_c23 :  std_logic_vector(35 downto 0);
signal expZm1adderX_c19 :  std_logic_vector(46 downto 0);
signal expZm1adderY_c23 :  std_logic_vector(46 downto 0);
signal expZm1_c24 :  std_logic_vector(46 downto 0);
signal expArounded_c20 :  std_logic_vector(45 downto 0);
signal lowerProduct_c26 :  std_logic_vector(47 downto 0);
signal extendedLowerProduct_c26 :  std_logic_vector(56 downto 0);
signal XSign_c15, XSign_c16, XSign_c17, XSign_c18 :  std_logic;
constant g: positive := 4;
constant wE: positive := 11;
constant wF: positive := 52;
constant wFIn: positive := 52;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_15 = '1' then
               XSign_c15 <= XSign;
            end if;
            if ce_16 = '1' then
               XSign_c16 <= XSign_c15;
            end if;
            if ce_17 = '1' then
               XSign_c17 <= XSign_c16;
            end if;
            if ce_18 = '1' then
               absK_c18 <= absK_c17;
               XSign_c18 <= XSign_c17;
            end if;
            if ce_19 = '1' then
            end if;
            if ce_20 = '1' then
            end if;
            if ce_21 = '1' then
            end if;
            if ce_22 = '1' then
            end if;
            if ce_23 = '1' then
            end if;
            if ce_24 = '1' then
            end if;
            if ce_25 = '1' then
            end if;
            if ce_26 = '1' then
            end if;
            if ce_27 = '1' then
            end if;
         end if;
      end process;
ufixX_c17 <= unsigned(ufixX_i);
   xMulIn_c17 <= ufixX_c17(65 downto 53); -- fix resize from (9, -56) to (9, -3)
   MulInvLog2: FixRealKCM_Freq300_uid1483
      port map ( clk  => clk,
                 X => std_logic_vector(xMulIn_c17),
                 R => absK_c17);
   minusAbsK_c18 <= (11 downto 0 => '0') - ('0' & absK_c18);
   K <= minusAbsK_c18 when  XSign_c18='1'   else ('0' & absK_c18);
   MulLog2: FixRealKCM_Freq300_uid1510
      port map ( clk  => clk,
                 ce_18 => ce_18,
                 X => absK_c17,
                 R => absKLog2_c18);
   subOp1_c17 <= std_logic_vector(ufixX_c17(55 downto 0)) when XSign_c17='0' else not (std_logic_vector(ufixX_c17(55 downto 0)));
   subOp2_c18 <= absKLog2_c18(55 downto 0) when XSign_c18='1' else not (absKLog2_c18(55 downto 0));
   theYAdder: IntAdder_56_Freq300_uid1523
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 Cin => '1',
                 X => subOp1_c17,
                 Y => subOp2_c18,
                 R => Y_c19);
   -- Now compute the exp of this fixed-point value
   A_c19 <= Y_c19(55 downto 46);
   Z_c19 <= Y_c19(45 downto 0);
   ExpATable: FixFunctionByTable_Freq300_uid1525
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 X => A_c19,
                 Y => expA_c20);
   Ztrunc_c19 <= Z_c19(45 downto 10);
   poly: FixFunctionByPiecewisePoly_Freq300_uid1534
      port map ( clk  => clk,
                 ce_20 => ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 X => Ztrunc_c19,
                 Y => expZmZm1_c23);
   -- Computing Z + (exp(Z)-1-Z)
   expZm1adderX_c19 <= '0' & Z_c19;
   expZm1adderY_c23 <= (10 downto 0 => '0') & expZmZm1_c23 ;
   Adder_expZm1: IntAdder_47_Freq300_uid2583
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 Cin => '0',
                 X => expZm1adderX_c19,
                 Y => expZm1adderY_c23,
                 R => expZm1_c24);
   -- Truncating expA to the same accuracy as expZm1
   expArounded_c20 <= expA_c20(56 downto 11);
   TheLowerProduct: IntMultiplier_46x47_48_Freq300_uid2585
      port map ( clk  => clk,
                 ce_21 => ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 X => expArounded_c20,
                 Y => expZm1_c24,
                 R => lowerProduct_c26);
   extendedLowerProduct_c26 <= ((56 downto 48 => '0') & lowerProduct_c26(47 downto 0));
   -- Final addition -- the product MSB bit weight is -k+2 = -8
   TheFinalAdder: IntAdder_57_Freq300_uid3177
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 Cin => '0',
                 X => expA_c20,
                 Y => extendedLowerProduct_c26,
                 R => expY);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_65_Freq300_uid3180
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq300_uid3180 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq300_uid3180 is
signal Rtmp_c27 :  std_logic_vector(64 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12, Cin_c13, Cin_c14, Cin_c15, Cin_c16, Cin_c17, Cin_c18, Cin_c19, Cin_c20, Cin_c21, Cin_c22, Cin_c23, Cin_c24, Cin_c25, Cin_c26, Cin_c27 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Cin_c12 <= Cin_c11;
            end if;
            if ce_13 = '1' then
               Cin_c13 <= Cin_c12;
            end if;
            if ce_14 = '1' then
               Cin_c14 <= Cin_c13;
            end if;
            if ce_15 = '1' then
               Cin_c15 <= Cin_c14;
            end if;
            if ce_16 = '1' then
               Cin_c16 <= Cin_c15;
            end if;
            if ce_17 = '1' then
               Cin_c17 <= Cin_c16;
            end if;
            if ce_18 = '1' then
               Cin_c18 <= Cin_c17;
            end if;
            if ce_19 = '1' then
               Cin_c19 <= Cin_c18;
            end if;
            if ce_20 = '1' then
               Cin_c20 <= Cin_c19;
            end if;
            if ce_21 = '1' then
               Cin_c21 <= Cin_c20;
            end if;
            if ce_22 = '1' then
               Cin_c22 <= Cin_c21;
            end if;
            if ce_23 = '1' then
               Cin_c23 <= Cin_c22;
            end if;
            if ce_24 = '1' then
               Cin_c24 <= Cin_c23;
            end if;
            if ce_25 = '1' then
               Cin_c25 <= Cin_c24;
            end if;
            if ce_26 = '1' then
               Cin_c26 <= Cin_c25;
            end if;
            if ce_27 = '1' then
               Cin_c27 <= Cin_c26;
            end if;
         end if;
      end process;
   Rtmp_c27 <= X + Y + Cin_c27;
   R <= Rtmp_c27;
end architecture;

--------------------------------------------------------------------------------
--                        FPExp_11_52_Freq300_uid1477
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPExp_11_52_Freq300_uid1477 is
    port (clk, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28 : in std_logic;
          X : in  std_logic_vector(11+67+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FPExp_11_52_Freq300_uid1477 is
   component LeftShifter68_by_max_65_Freq300_uid1479 is
      port ( clk, ce_15, ce_16, ce_17 : in std_logic;
             X : in  std_logic_vector(67 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(132 downto 0)   );
   end component;

   component Exp_11_52_Freq300_uid1481 is
      port ( clk, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27 : in std_logic;
             ufixX_i : in  std_logic_vector(65 downto 0);
             XSign : in  std_logic;
             expY : out  std_logic_vector(56 downto 0);
             K : out  std_logic_vector(11 downto 0)   );
   end component;

   component IntAdder_65_Freq300_uid3180 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal Xexn_c14, Xexn_c15, Xexn_c16, Xexn_c17, Xexn_c18, Xexn_c19, Xexn_c20, Xexn_c21, Xexn_c22, Xexn_c23, Xexn_c24, Xexn_c25, Xexn_c26, Xexn_c27, Xexn_c28 :  std_logic_vector(1 downto 0);
signal XSign_c14, XSign_c15, XSign_c16, XSign_c17, XSign_c18, XSign_c19, XSign_c20, XSign_c21, XSign_c22, XSign_c23, XSign_c24, XSign_c25, XSign_c26, XSign_c27, XSign_c28 :  std_logic;
signal XexpField_c14, XexpField_c15 :  std_logic_vector(10 downto 0);
signal Xfrac_c14 :  unsigned(-1+67 downto 0);
signal e0_c0, e0_c1, e0_c2, e0_c3, e0_c4, e0_c5, e0_c6, e0_c7, e0_c8, e0_c9, e0_c10, e0_c11, e0_c12, e0_c13, e0_c14, e0_c15 :  std_logic_vector(12 downto 0);
signal shiftVal_c15 :  std_logic_vector(12 downto 0);
signal resultWillBeOne_c15, resultWillBeOne_c16, resultWillBeOne_c17 :  std_logic;
signal mXu_c14 :  unsigned(0+67 downto 0);
signal maxShift_c0, maxShift_c1, maxShift_c2, maxShift_c3, maxShift_c4, maxShift_c5, maxShift_c6, maxShift_c7, maxShift_c8, maxShift_c9, maxShift_c10, maxShift_c11, maxShift_c12, maxShift_c13, maxShift_c14, maxShift_c15 :  std_logic_vector(11 downto 0);
signal overflow0_c15 :  std_logic;
signal shiftValIn_c15 :  std_logic_vector(6 downto 0);
signal fixX0_c17 :  std_logic_vector(132 downto 0);
signal ufixX_c17 :  unsigned(9+56 downto 0);
signal expY_c27 :  std_logic_vector(56 downto 0);
signal K_c18, K_c19, K_c20, K_c21, K_c22, K_c23, K_c24, K_c25, K_c26, K_c27 :  std_logic_vector(11 downto 0);
signal needNoNorm_c27 :  std_logic;
signal preRoundBiasSig_c27 :  std_logic_vector(64 downto 0);
signal roundBit_c27 :  std_logic;
signal roundNormAddend_c27 :  std_logic_vector(64 downto 0);
signal roundedExpSigRes_c27, roundedExpSigRes_c28 :  std_logic_vector(64 downto 0);
signal roundedExpSig_c28 :  std_logic_vector(64 downto 0);
signal ofl1_c15, ofl1_c16, ofl1_c17, ofl1_c18, ofl1_c19, ofl1_c20, ofl1_c21, ofl1_c22, ofl1_c23, ofl1_c24, ofl1_c25, ofl1_c26, ofl1_c27, ofl1_c28 :  std_logic;
signal ofl2_c28 :  std_logic;
signal ofl3_c14, ofl3_c15, ofl3_c16, ofl3_c17, ofl3_c18, ofl3_c19, ofl3_c20, ofl3_c21, ofl3_c22, ofl3_c23, ofl3_c24, ofl3_c25, ofl3_c26, ofl3_c27, ofl3_c28 :  std_logic;
signal ofl_c28 :  std_logic;
signal ufl1_c28 :  std_logic;
signal ufl2_c14, ufl2_c15, ufl2_c16, ufl2_c17, ufl2_c18, ufl2_c19, ufl2_c20, ufl2_c21, ufl2_c22, ufl2_c23, ufl2_c24, ufl2_c25, ufl2_c26, ufl2_c27, ufl2_c28 :  std_logic;
signal ufl3_c15, ufl3_c16, ufl3_c17, ufl3_c18, ufl3_c19, ufl3_c20, ufl3_c21, ufl3_c22, ufl3_c23, ufl3_c24, ufl3_c25, ufl3_c26, ufl3_c27, ufl3_c28 :  std_logic;
signal ufl_c28 :  std_logic;
signal Rexn_c28 :  std_logic_vector(1 downto 0);
constant g: positive := 4;
constant wE: positive := 11;
constant wF: positive := 52;
constant wFIn: positive := 67;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_15 = '1' then
               Xexn_c15 <= Xexn_c14;
               XSign_c15 <= XSign_c14;
               XexpField_c15 <= XexpField_c14;
               e0_c15 <= e0_c14;
               maxShift_c15 <= maxShift_c14;
               ofl3_c15 <= ofl3_c14;
               ufl2_c15 <= ufl2_c14;
            end if;
            if ce_16 = '1' then
               Xexn_c16 <= Xexn_c15;
               XSign_c16 <= XSign_c15;
               resultWillBeOne_c16 <= resultWillBeOne_c15;
               ofl1_c16 <= ofl1_c15;
               ofl3_c16 <= ofl3_c15;
               ufl2_c16 <= ufl2_c15;
               ufl3_c16 <= ufl3_c15;
            end if;
            if ce_17 = '1' then
               Xexn_c17 <= Xexn_c16;
               XSign_c17 <= XSign_c16;
               resultWillBeOne_c17 <= resultWillBeOne_c16;
               ofl1_c17 <= ofl1_c16;
               ofl3_c17 <= ofl3_c16;
               ufl2_c17 <= ufl2_c16;
               ufl3_c17 <= ufl3_c16;
            end if;
            if ce_18 = '1' then
               Xexn_c18 <= Xexn_c17;
               XSign_c18 <= XSign_c17;
               ofl1_c18 <= ofl1_c17;
               ofl3_c18 <= ofl3_c17;
               ufl2_c18 <= ufl2_c17;
               ufl3_c18 <= ufl3_c17;
            end if;
            if ce_19 = '1' then
               Xexn_c19 <= Xexn_c18;
               XSign_c19 <= XSign_c18;
               K_c19 <= K_c18;
               ofl1_c19 <= ofl1_c18;
               ofl3_c19 <= ofl3_c18;
               ufl2_c19 <= ufl2_c18;
               ufl3_c19 <= ufl3_c18;
            end if;
            if ce_20 = '1' then
               Xexn_c20 <= Xexn_c19;
               XSign_c20 <= XSign_c19;
               K_c20 <= K_c19;
               ofl1_c20 <= ofl1_c19;
               ofl3_c20 <= ofl3_c19;
               ufl2_c20 <= ufl2_c19;
               ufl3_c20 <= ufl3_c19;
            end if;
            if ce_21 = '1' then
               Xexn_c21 <= Xexn_c20;
               XSign_c21 <= XSign_c20;
               K_c21 <= K_c20;
               ofl1_c21 <= ofl1_c20;
               ofl3_c21 <= ofl3_c20;
               ufl2_c21 <= ufl2_c20;
               ufl3_c21 <= ufl3_c20;
            end if;
            if ce_22 = '1' then
               Xexn_c22 <= Xexn_c21;
               XSign_c22 <= XSign_c21;
               K_c22 <= K_c21;
               ofl1_c22 <= ofl1_c21;
               ofl3_c22 <= ofl3_c21;
               ufl2_c22 <= ufl2_c21;
               ufl3_c22 <= ufl3_c21;
            end if;
            if ce_23 = '1' then
               Xexn_c23 <= Xexn_c22;
               XSign_c23 <= XSign_c22;
               K_c23 <= K_c22;
               ofl1_c23 <= ofl1_c22;
               ofl3_c23 <= ofl3_c22;
               ufl2_c23 <= ufl2_c22;
               ufl3_c23 <= ufl3_c22;
            end if;
            if ce_24 = '1' then
               Xexn_c24 <= Xexn_c23;
               XSign_c24 <= XSign_c23;
               K_c24 <= K_c23;
               ofl1_c24 <= ofl1_c23;
               ofl3_c24 <= ofl3_c23;
               ufl2_c24 <= ufl2_c23;
               ufl3_c24 <= ufl3_c23;
            end if;
            if ce_25 = '1' then
               Xexn_c25 <= Xexn_c24;
               XSign_c25 <= XSign_c24;
               K_c25 <= K_c24;
               ofl1_c25 <= ofl1_c24;
               ofl3_c25 <= ofl3_c24;
               ufl2_c25 <= ufl2_c24;
               ufl3_c25 <= ufl3_c24;
            end if;
            if ce_26 = '1' then
               Xexn_c26 <= Xexn_c25;
               XSign_c26 <= XSign_c25;
               K_c26 <= K_c25;
               ofl1_c26 <= ofl1_c25;
               ofl3_c26 <= ofl3_c25;
               ufl2_c26 <= ufl2_c25;
               ufl3_c26 <= ufl3_c25;
            end if;
            if ce_27 = '1' then
               Xexn_c27 <= Xexn_c26;
               XSign_c27 <= XSign_c26;
               K_c27 <= K_c26;
               ofl1_c27 <= ofl1_c26;
               ofl3_c27 <= ofl3_c26;
               ufl2_c27 <= ufl2_c26;
               ufl3_c27 <= ufl3_c26;
            end if;
            if ce_28 = '1' then
               Xexn_c28 <= Xexn_c27;
               XSign_c28 <= XSign_c27;
               roundedExpSigRes_c28 <= roundedExpSigRes_c27;
               ofl1_c28 <= ofl1_c27;
               ofl3_c28 <= ofl3_c27;
               ufl2_c28 <= ufl2_c27;
               ufl3_c28 <= ufl3_c27;
            end if;
         end if;
      end process;
   Xexn_c14 <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign_c14 <= X(wE+wFIn);
   XexpField_c14 <= X(wE+wFIn-1 downto wFIn);
   Xfrac_c14 <= unsigned(X(wFIn-1 downto 0));
   e0_c0 <= conv_std_logic_vector(967, wE+2);  -- bias - (wF+g)
   shiftVal_c15 <= ("00" & XexpField_c15) - e0_c15; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne_c15 <= shiftVal_c15(wE+1);
   --  mantissa with implicit bit
   mXu_c14 <= "1" & Xfrac_c14;
   -- Partial overflow detection
   maxShift_c0 <= conv_std_logic_vector(65, wE+1);  -- wE-2 + wF+g
   overflow0_c15 <= not shiftVal_c15(wE+1) when shiftVal_c15(wE downto 0) > maxShift_c15 else '0';
   shiftValIn_c15 <= shiftVal_c15(6 downto 0);
   mantissa_shift: LeftShifter68_by_max_65_Freq300_uid1479
      port map ( clk  => clk,
                 ce_15 => ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 S => shiftValIn_c15,
                 X => std_logic_vector(mXu_c14),
                 R => fixX0_c17);
   ufixX_c17 <=  unsigned(fixX0_c17(132 downto 67)) when resultWillBeOne_c17='0' else "000000000000000000000000000000000000000000000000000000000000000000";
   exp_helper: Exp_11_52_Freq300_uid1481
      port map ( clk  => clk,
                 ce_15 => ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 XSign => XSign_c14,
                 ufixX_i => std_logic_vector(ufixX_c17),
                 K => K_c18,
                 expY => expY_c27);
   needNoNorm_c27 <= expY_c27(56);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig_c27 <= conv_std_logic_vector(1023, wE+2)  & expY_c27(55 downto 4) when needNoNorm_c27 = '1'
      else conv_std_logic_vector(1022, wE+2)  & expY_c27(54 downto 3) ;
   roundBit_c27 <= expY_c27(3)  when needNoNorm_c27 = '1'    else expY_c27(2) ;
   roundNormAddend_c27 <= K_c27(11) & K_c27 & (51 downto 1 => '0') & roundBit_c27;
   roundedExpSigOperandAdder: IntAdder_65_Freq300_uid3180
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 Cin => '0',
                 X => preRoundBiasSig_c27,
                 Y => roundNormAddend_c27,
                 R => roundedExpSigRes_c27);
   roundedExpSig_c28 <= roundedExpSigRes_c28 when Xexn_c28="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1_c15 <= not XSign_c15 and overflow0_c15 and (not Xexn_c15(1) and Xexn_c15(0)); -- input positive, normal,  very large
   ofl2_c28 <= not XSign_c28 and (roundedExpSig_c28(wE+wF) and not roundedExpSig_c28(wE+wF+1)) and (not Xexn_c28(1) and Xexn_c28(0)); -- input positive, normal, overflowed
   ofl3_c14 <= not XSign_c14 and Xexn_c14(1) and not Xexn_c14(0);  -- input was -infty
   ofl_c28 <= ofl1_c28 or ofl2_c28 or ofl3_c28;
   ufl1_c28 <= (roundedExpSig_c28(wE+wF) and roundedExpSig_c28(wE+wF+1))  and (not Xexn_c28(1) and Xexn_c28(0)); -- input normal
   ufl2_c14 <= XSign_c14 and Xexn_c14(1) and not Xexn_c14(0);  -- input was -infty
   ufl3_c15 <= XSign_c15 and overflow0_c15  and (not Xexn_c15(1) and Xexn_c15(0)); -- input negative, normal,  very large
   ufl_c28 <= ufl1_c28 or ufl2_c28 or ufl3_c28;
   Rexn_c28 <= "11" when Xexn_c28 = "11"
      else "10" when ofl_c28='1'
      else "00" when ufl_c28='1'
      else "01";
   R <= Rexn_c28 & '0' & roundedExpSig_c28(62 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointPower
--                         (FPPow_11_52_Freq300_uid2)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointPower is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointPower is
   component IntAdder_64_Freq300_uid5 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(63 downto 0);
             Y : in  std_logic_vector(63 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(63 downto 0)   );
   end component;

   component LZC_52_Freq300_uid7 is
      port ( clk, ce_1 : in std_logic;
             I : in  std_logic_vector(51 downto 0);
             O : out  std_logic_vector(5 downto 0)   );
   end component;

   component FPLogIterative_11_66_0_300_Freq300_uid9 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(11+66+2 downto 0);
             R : out  std_logic_vector(11+66+2 downto 0)   );
   end component;

   component FPMult_11_66_uid81_Freq300_uid82 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14 : in std_logic;
             X : in  std_logic_vector(11+66+2 downto 0);
             Y : in  std_logic_vector(11+52+2 downto 0);
             R : out  std_logic_vector(11+67+2 downto 0)   );
   end component;

   component FPExp_11_52_Freq300_uid1477 is
      port ( clk, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28 : in std_logic;
             X : in  std_logic_vector(11+67+2 downto 0);
             R : out  std_logic_vector(11+52+2 downto 0)   );
   end component;

signal flagsX_c0 :  std_logic_vector(1 downto 0);
signal signX_c0, signX_c1, signX_c2 :  std_logic;
signal expFieldX_c0 :  std_logic_vector(10 downto 0);
signal fracX_c0 :  std_logic_vector(51 downto 0);
signal flagsY_c0 :  std_logic_vector(1 downto 0);
signal signY_c0, signY_c1, signY_c2 :  std_logic;
signal expFieldY_c0 :  std_logic_vector(10 downto 0);
signal fracY_c0 :  std_logic_vector(51 downto 0);
signal zeroX_c0, zeroX_c1, zeroX_c2 :  std_logic;
signal zeroY_c0, zeroY_c1, zeroY_c2 :  std_logic;
signal normalX_c0, normalX_c1, normalX_c2 :  std_logic;
signal normalY_c0, normalY_c1, normalY_c2 :  std_logic;
signal infX_c0, infX_c1, infX_c2 :  std_logic;
signal infY_c0, infY_c1, infY_c2 :  std_logic;
signal s_nan_in_c0, s_nan_in_c1, s_nan_in_c2 :  std_logic;
signal OneExpFrac_c0 :  std_logic_vector(62 downto 0);
signal ExpFracX_c0 :  std_logic_vector(63 downto 0);
signal OneExpFracCompl_c0 :  std_logic_vector(63 downto 0);
signal cmpXOneRes_c0 :  std_logic_vector(63 downto 0);
signal XisOneAndNormal_c0 :  std_logic;
signal absXgtOneAndNormal_c0, absXgtOneAndNormal_c1, absXgtOneAndNormal_c2 :  std_logic;
signal absXltOneAndNormal_c0, absXltOneAndNormal_c1, absXltOneAndNormal_c2 :  std_logic;
signal fracYreverted_c0 :  std_logic_vector(51 downto 0);
signal Z_rightY_c1 :  std_logic_vector(5 downto 0);
signal WeightLSBYpre_c0, WeightLSBYpre_c1 :  std_logic_vector(11 downto 0);
signal WeightLSBY_c1, WeightLSBY_c2 :  std_logic_vector(11 downto 0);
signal oddIntY_c2 :  std_logic;
signal evenIntY_c2 :  std_logic;
signal notIntNormalY_c2 :  std_logic;
signal RisInfSpecialCase_c2, RisInfSpecialCase_c3, RisInfSpecialCase_c4, RisInfSpecialCase_c5, RisInfSpecialCase_c6, RisInfSpecialCase_c7, RisInfSpecialCase_c8, RisInfSpecialCase_c9, RisInfSpecialCase_c10, RisInfSpecialCase_c11, RisInfSpecialCase_c12, RisInfSpecialCase_c13, RisInfSpecialCase_c14, RisInfSpecialCase_c15, RisInfSpecialCase_c16, RisInfSpecialCase_c17, RisInfSpecialCase_c18, RisInfSpecialCase_c19, RisInfSpecialCase_c20, RisInfSpecialCase_c21, RisInfSpecialCase_c22, RisInfSpecialCase_c23, RisInfSpecialCase_c24, RisInfSpecialCase_c25, RisInfSpecialCase_c26, RisInfSpecialCase_c27, RisInfSpecialCase_c28 :  std_logic;
signal RisZeroSpecialCase_c2, RisZeroSpecialCase_c3, RisZeroSpecialCase_c4, RisZeroSpecialCase_c5, RisZeroSpecialCase_c6, RisZeroSpecialCase_c7, RisZeroSpecialCase_c8, RisZeroSpecialCase_c9, RisZeroSpecialCase_c10, RisZeroSpecialCase_c11, RisZeroSpecialCase_c12, RisZeroSpecialCase_c13, RisZeroSpecialCase_c14, RisZeroSpecialCase_c15, RisZeroSpecialCase_c16, RisZeroSpecialCase_c17, RisZeroSpecialCase_c18, RisZeroSpecialCase_c19, RisZeroSpecialCase_c20, RisZeroSpecialCase_c21, RisZeroSpecialCase_c22, RisZeroSpecialCase_c23, RisZeroSpecialCase_c24, RisZeroSpecialCase_c25, RisZeroSpecialCase_c26, RisZeroSpecialCase_c27, RisZeroSpecialCase_c28 :  std_logic;
signal RisOne_c0, RisOne_c1, RisOne_c2, RisOne_c3, RisOne_c4, RisOne_c5, RisOne_c6, RisOne_c7, RisOne_c8, RisOne_c9, RisOne_c10, RisOne_c11, RisOne_c12, RisOne_c13, RisOne_c14, RisOne_c15, RisOne_c16, RisOne_c17, RisOne_c18, RisOne_c19, RisOne_c20, RisOne_c21, RisOne_c22, RisOne_c23, RisOne_c24, RisOne_c25, RisOne_c26, RisOne_c27, RisOne_c28 :  std_logic;
signal RisNaN_c2, RisNaN_c3, RisNaN_c4, RisNaN_c5, RisNaN_c6, RisNaN_c7, RisNaN_c8, RisNaN_c9, RisNaN_c10, RisNaN_c11, RisNaN_c12, RisNaN_c13, RisNaN_c14, RisNaN_c15, RisNaN_c16, RisNaN_c17, RisNaN_c18, RisNaN_c19, RisNaN_c20, RisNaN_c21, RisNaN_c22, RisNaN_c23, RisNaN_c24, RisNaN_c25, RisNaN_c26, RisNaN_c27, RisNaN_c28 :  std_logic;
signal signR_c2, signR_c3, signR_c4, signR_c5, signR_c6, signR_c7, signR_c8, signR_c9, signR_c10, signR_c11, signR_c12, signR_c13, signR_c14, signR_c15, signR_c16, signR_c17, signR_c18, signR_c19, signR_c20, signR_c21, signR_c22, signR_c23, signR_c24, signR_c25, signR_c26, signR_c27, signR_c28 :  std_logic;
signal logIn_c0 :  std_logic_vector(79 downto 0);
signal lnX_c11 :  std_logic_vector(11+66+2 downto 0);
signal P_c14 :  std_logic_vector(11+67+2 downto 0);
signal E_c28 :  std_logic_vector(11+52+2 downto 0);
signal flagsE_c28 :  std_logic_vector(1 downto 0);
signal RisZeroFromExp_c28 :  std_logic;
signal RisZero_c28 :  std_logic;
signal RisInfFromExp_c28 :  std_logic;
signal RisInf_c28 :  std_logic;
signal flagR_c28 :  std_logic_vector(1 downto 0);
signal R_expfrac_c28 :  std_logic_vector(62 downto 0);
constant wE: positive := 11;
constant wF: positive := 52;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               signX_c1 <= signX_c0;
               signY_c1 <= signY_c0;
               zeroX_c1 <= zeroX_c0;
               zeroY_c1 <= zeroY_c0;
               normalX_c1 <= normalX_c0;
               normalY_c1 <= normalY_c0;
               infX_c1 <= infX_c0;
               infY_c1 <= infY_c0;
               s_nan_in_c1 <= s_nan_in_c0;
               absXgtOneAndNormal_c1 <= absXgtOneAndNormal_c0;
               absXltOneAndNormal_c1 <= absXltOneAndNormal_c0;
               WeightLSBYpre_c1 <= WeightLSBYpre_c0;
               RisOne_c1 <= RisOne_c0;
            end if;
            if ce_2 = '1' then
               signX_c2 <= signX_c1;
               signY_c2 <= signY_c1;
               zeroX_c2 <= zeroX_c1;
               zeroY_c2 <= zeroY_c1;
               normalX_c2 <= normalX_c1;
               normalY_c2 <= normalY_c1;
               infX_c2 <= infX_c1;
               infY_c2 <= infY_c1;
               s_nan_in_c2 <= s_nan_in_c1;
               absXgtOneAndNormal_c2 <= absXgtOneAndNormal_c1;
               absXltOneAndNormal_c2 <= absXltOneAndNormal_c1;
               WeightLSBY_c2 <= WeightLSBY_c1;
               RisOne_c2 <= RisOne_c1;
            end if;
            if ce_3 = '1' then
               RisInfSpecialCase_c3 <= RisInfSpecialCase_c2;
               RisZeroSpecialCase_c3 <= RisZeroSpecialCase_c2;
               RisOne_c3 <= RisOne_c2;
               RisNaN_c3 <= RisNaN_c2;
               signR_c3 <= signR_c2;
            end if;
            if ce_4 = '1' then
               RisInfSpecialCase_c4 <= RisInfSpecialCase_c3;
               RisZeroSpecialCase_c4 <= RisZeroSpecialCase_c3;
               RisOne_c4 <= RisOne_c3;
               RisNaN_c4 <= RisNaN_c3;
               signR_c4 <= signR_c3;
            end if;
            if ce_5 = '1' then
               RisInfSpecialCase_c5 <= RisInfSpecialCase_c4;
               RisZeroSpecialCase_c5 <= RisZeroSpecialCase_c4;
               RisOne_c5 <= RisOne_c4;
               RisNaN_c5 <= RisNaN_c4;
               signR_c5 <= signR_c4;
            end if;
            if ce_6 = '1' then
               RisInfSpecialCase_c6 <= RisInfSpecialCase_c5;
               RisZeroSpecialCase_c6 <= RisZeroSpecialCase_c5;
               RisOne_c6 <= RisOne_c5;
               RisNaN_c6 <= RisNaN_c5;
               signR_c6 <= signR_c5;
            end if;
            if ce_7 = '1' then
               RisInfSpecialCase_c7 <= RisInfSpecialCase_c6;
               RisZeroSpecialCase_c7 <= RisZeroSpecialCase_c6;
               RisOne_c7 <= RisOne_c6;
               RisNaN_c7 <= RisNaN_c6;
               signR_c7 <= signR_c6;
            end if;
            if ce_8 = '1' then
               RisInfSpecialCase_c8 <= RisInfSpecialCase_c7;
               RisZeroSpecialCase_c8 <= RisZeroSpecialCase_c7;
               RisOne_c8 <= RisOne_c7;
               RisNaN_c8 <= RisNaN_c7;
               signR_c8 <= signR_c7;
            end if;
            if ce_9 = '1' then
               RisInfSpecialCase_c9 <= RisInfSpecialCase_c8;
               RisZeroSpecialCase_c9 <= RisZeroSpecialCase_c8;
               RisOne_c9 <= RisOne_c8;
               RisNaN_c9 <= RisNaN_c8;
               signR_c9 <= signR_c8;
            end if;
            if ce_10 = '1' then
               RisInfSpecialCase_c10 <= RisInfSpecialCase_c9;
               RisZeroSpecialCase_c10 <= RisZeroSpecialCase_c9;
               RisOne_c10 <= RisOne_c9;
               RisNaN_c10 <= RisNaN_c9;
               signR_c10 <= signR_c9;
            end if;
            if ce_11 = '1' then
               RisInfSpecialCase_c11 <= RisInfSpecialCase_c10;
               RisZeroSpecialCase_c11 <= RisZeroSpecialCase_c10;
               RisOne_c11 <= RisOne_c10;
               RisNaN_c11 <= RisNaN_c10;
               signR_c11 <= signR_c10;
            end if;
            if ce_12 = '1' then
               RisInfSpecialCase_c12 <= RisInfSpecialCase_c11;
               RisZeroSpecialCase_c12 <= RisZeroSpecialCase_c11;
               RisOne_c12 <= RisOne_c11;
               RisNaN_c12 <= RisNaN_c11;
               signR_c12 <= signR_c11;
            end if;
            if ce_13 = '1' then
               RisInfSpecialCase_c13 <= RisInfSpecialCase_c12;
               RisZeroSpecialCase_c13 <= RisZeroSpecialCase_c12;
               RisOne_c13 <= RisOne_c12;
               RisNaN_c13 <= RisNaN_c12;
               signR_c13 <= signR_c12;
            end if;
            if ce_14 = '1' then
               RisInfSpecialCase_c14 <= RisInfSpecialCase_c13;
               RisZeroSpecialCase_c14 <= RisZeroSpecialCase_c13;
               RisOne_c14 <= RisOne_c13;
               RisNaN_c14 <= RisNaN_c13;
               signR_c14 <= signR_c13;
            end if;
            if ce_15 = '1' then
               RisInfSpecialCase_c15 <= RisInfSpecialCase_c14;
               RisZeroSpecialCase_c15 <= RisZeroSpecialCase_c14;
               RisOne_c15 <= RisOne_c14;
               RisNaN_c15 <= RisNaN_c14;
               signR_c15 <= signR_c14;
            end if;
            if ce_16 = '1' then
               RisInfSpecialCase_c16 <= RisInfSpecialCase_c15;
               RisZeroSpecialCase_c16 <= RisZeroSpecialCase_c15;
               RisOne_c16 <= RisOne_c15;
               RisNaN_c16 <= RisNaN_c15;
               signR_c16 <= signR_c15;
            end if;
            if ce_17 = '1' then
               RisInfSpecialCase_c17 <= RisInfSpecialCase_c16;
               RisZeroSpecialCase_c17 <= RisZeroSpecialCase_c16;
               RisOne_c17 <= RisOne_c16;
               RisNaN_c17 <= RisNaN_c16;
               signR_c17 <= signR_c16;
            end if;
            if ce_18 = '1' then
               RisInfSpecialCase_c18 <= RisInfSpecialCase_c17;
               RisZeroSpecialCase_c18 <= RisZeroSpecialCase_c17;
               RisOne_c18 <= RisOne_c17;
               RisNaN_c18 <= RisNaN_c17;
               signR_c18 <= signR_c17;
            end if;
            if ce_19 = '1' then
               RisInfSpecialCase_c19 <= RisInfSpecialCase_c18;
               RisZeroSpecialCase_c19 <= RisZeroSpecialCase_c18;
               RisOne_c19 <= RisOne_c18;
               RisNaN_c19 <= RisNaN_c18;
               signR_c19 <= signR_c18;
            end if;
            if ce_20 = '1' then
               RisInfSpecialCase_c20 <= RisInfSpecialCase_c19;
               RisZeroSpecialCase_c20 <= RisZeroSpecialCase_c19;
               RisOne_c20 <= RisOne_c19;
               RisNaN_c20 <= RisNaN_c19;
               signR_c20 <= signR_c19;
            end if;
            if ce_21 = '1' then
               RisInfSpecialCase_c21 <= RisInfSpecialCase_c20;
               RisZeroSpecialCase_c21 <= RisZeroSpecialCase_c20;
               RisOne_c21 <= RisOne_c20;
               RisNaN_c21 <= RisNaN_c20;
               signR_c21 <= signR_c20;
            end if;
            if ce_22 = '1' then
               RisInfSpecialCase_c22 <= RisInfSpecialCase_c21;
               RisZeroSpecialCase_c22 <= RisZeroSpecialCase_c21;
               RisOne_c22 <= RisOne_c21;
               RisNaN_c22 <= RisNaN_c21;
               signR_c22 <= signR_c21;
            end if;
            if ce_23 = '1' then
               RisInfSpecialCase_c23 <= RisInfSpecialCase_c22;
               RisZeroSpecialCase_c23 <= RisZeroSpecialCase_c22;
               RisOne_c23 <= RisOne_c22;
               RisNaN_c23 <= RisNaN_c22;
               signR_c23 <= signR_c22;
            end if;
            if ce_24 = '1' then
               RisInfSpecialCase_c24 <= RisInfSpecialCase_c23;
               RisZeroSpecialCase_c24 <= RisZeroSpecialCase_c23;
               RisOne_c24 <= RisOne_c23;
               RisNaN_c24 <= RisNaN_c23;
               signR_c24 <= signR_c23;
            end if;
            if ce_25 = '1' then
               RisInfSpecialCase_c25 <= RisInfSpecialCase_c24;
               RisZeroSpecialCase_c25 <= RisZeroSpecialCase_c24;
               RisOne_c25 <= RisOne_c24;
               RisNaN_c25 <= RisNaN_c24;
               signR_c25 <= signR_c24;
            end if;
            if ce_26 = '1' then
               RisInfSpecialCase_c26 <= RisInfSpecialCase_c25;
               RisZeroSpecialCase_c26 <= RisZeroSpecialCase_c25;
               RisOne_c26 <= RisOne_c25;
               RisNaN_c26 <= RisNaN_c25;
               signR_c26 <= signR_c25;
            end if;
            if ce_27 = '1' then
               RisInfSpecialCase_c27 <= RisInfSpecialCase_c26;
               RisZeroSpecialCase_c27 <= RisZeroSpecialCase_c26;
               RisOne_c27 <= RisOne_c26;
               RisNaN_c27 <= RisNaN_c26;
               signR_c27 <= signR_c26;
            end if;
            if ce_28 = '1' then
               RisInfSpecialCase_c28 <= RisInfSpecialCase_c27;
               RisZeroSpecialCase_c28 <= RisZeroSpecialCase_c27;
               RisOne_c28 <= RisOne_c27;
               RisNaN_c28 <= RisNaN_c27;
               signR_c28 <= signR_c27;
            end if;
         end if;
      end process;
   flagsX_c0 <= X(wE+wF+2 downto wE+wF+1);
   signX_c0 <= X(wE+wF);
   expFieldX_c0 <= X(wE+wF-1 downto wF);
   fracX_c0 <= X(wF-1 downto 0);
   flagsY_c0 <= Y(wE+wF+2 downto wE+wF+1);
   signY_c0 <= Y(wE+wF);
   expFieldY_c0 <= Y(wE+wF-1 downto wF);
   fracY_c0 <= Y(wF-1 downto 0);
-- Inputs analysis  --
-- zero inputs--
   zeroX_c0 <= '1' when flagsX_c0="00" else '0';
   zeroY_c0 <= '1' when flagsY_c0="00" else '0';
-- normal inputs--
   normalX_c0 <= '1' when flagsX_c0="01" else '0';
   normalY_c0 <= '1' when flagsY_c0="01" else '0';
-- inf input --
   infX_c0 <= '1' when flagsX_c0="10" else '0';
   infY_c0 <= '1' when flagsY_c0="10" else '0';
-- NaN inputs  --
   s_nan_in_c0 <= '1' when flagsX_c0="11" or flagsY_c0="11" else '0';
-- Comparison of X to 1   --
   OneExpFrac_c0 <=  "0" & (9 downto 0 => '1') & (51 downto 0 => '0');
   ExpFracX_c0<= "0" & expFieldX_c0 & fracX_c0;
   OneExpFracCompl_c0<=  "1" & (not OneExpFrac_c0);
   cmpXOne: IntAdder_64_Freq300_uid5
      port map ( clk  => clk,
                 Cin => '1',
                 X => ExpFracX_c0,
                 Y => OneExpFracCompl_c0,
                 R => cmpXOneRes_c0);
   XisOneAndNormal_c0 <= '1' when X = ("010" & OneExpFrac_c0) else '0';
   absXgtOneAndNormal_c0 <= normalX_c0 and (not XisOneAndNormal_c0) and (not cmpXOneRes_c0(63));
   absXltOneAndNormal_c0 <= normalX_c0 and cmpXOneRes_c0(63);
   fracYreverted_c0 <= fracY_c0(0)&fracY_c0(1)&fracY_c0(2)&fracY_c0(3)&fracY_c0(4)&fracY_c0(5)&fracY_c0(6)&fracY_c0(7)&fracY_c0(8)&fracY_c0(9)&fracY_c0(10)&fracY_c0(11)&fracY_c0(12)&fracY_c0(13)&fracY_c0(14)&fracY_c0(15)&fracY_c0(16)&fracY_c0(17)&fracY_c0(18)&fracY_c0(19)&fracY_c0(20)&fracY_c0(21)&fracY_c0(22)&fracY_c0(23)&fracY_c0(24)&fracY_c0(25)&fracY_c0(26)&fracY_c0(27)&fracY_c0(28)&fracY_c0(29)&fracY_c0(30)&fracY_c0(31)&fracY_c0(32)&fracY_c0(33)&fracY_c0(34)&fracY_c0(35)&fracY_c0(36)&fracY_c0(37)&fracY_c0(38)&fracY_c0(39)&fracY_c0(40)&fracY_c0(41)&fracY_c0(42)&fracY_c0(43)&fracY_c0(44)&fracY_c0(45)&fracY_c0(46)&fracY_c0(47)&fracY_c0(48)&fracY_c0(49)&fracY_c0(50)&fracY_c0(51);
   FPPow_11_52_Freq300_uid2right1counter: LZC_52_Freq300_uid7
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 I => fracYreverted_c0,
                 O => Z_rightY_c1);
-- compute the weight of the less significant one of the mantissa
   WeightLSBYpre_c0 <= ('0' & expFieldY_c0)- CONV_STD_LOGIC_VECTOR(1075,12);
   WeightLSBY_c1 <= WeightLSBYpre_c1 + Z_rightY_c1;
   oddIntY_c2 <= normalY_c2 when WeightLSBY_c2 = CONV_STD_LOGIC_VECTOR(0, 12) else '0'; -- LSB has null weight
   evenIntY_c2 <= normalY_c2 when WeightLSBY_c2(wE)='0' and oddIntY_c2='0' else '0'; --LSB has strictly positive weight 
   notIntNormalY_c2 <= normalY_c2 when WeightLSBY_c2(wE)='1' else '0'; -- LSB has negative weight

-- Pow Exceptions  --
   RisInfSpecialCase_c2  <= 
         (zeroX_c2  and  (oddIntY_c2 or evenIntY_c2)  and signY_c2)  -- (+/- 0) ^ (negative int y)
      or (zeroX_c2 and infY_c2 and signY_c2)                      -- (+/- 0) ^ (-inf)
      or (absXgtOneAndNormal_c2   and  infY_c2  and not signY_c2) -- (|x|>1) ^ (+inf)
      or (absXltOneAndNormal_c2   and  infY_c2  and signY_c2)     -- (|x|<1) ^ (-inf)
      or (infX_c2 and  normalY_c2  and not signY_c2) ;            -- (inf) ^ (y>0)
   RisZeroSpecialCase_c2 <= 
         (zeroX_c2 and  (oddIntY_c2 or evenIntY_c2)  and not signY_c2)  -- (+/- 0) ^ (positive int y)
      or (zeroX_c2 and  infY_c2  and not signY_c2)                   -- (+/- 0) ^ (+inf)
      or (absXltOneAndNormal_c2   and  infY_c2  and not signY_c2)    -- (|x|<1) ^ (+inf)
      or (absXgtOneAndNormal_c2   and  infY_c2  and signY_c2)        -- (|x|>1) ^ (-inf)
      or (infX_c2 and  normalY_c2  and signY_c2) ;                   -- (inf) ^ (y<0)
   RisOne_c0 <= 
         zeroY_c0                                          -- x^0 = 1 without exception
      or (XisOneAndNormal_c0 and signX_c0 and infY_c0)           -- (-1) ^ (-/-inf)
      or (XisOneAndNormal_c0  and not signX_c0);              -- (+1) ^ (whatever)
   RisNaN_c2 <= (s_nan_in_c2 and not zeroY_c2) or (normalX_c2 and signX_c2 and notIntNormalY_c2);
   signR_c2 <= signX_c2 and (oddIntY_c2);
   logIn_c0 <= flagsX_c0 & "0" & expFieldX_c0 & fracX_c0 & (13 downto 0 => '0') ;
   FPPow_11_52_Freq300_uid2log: FPLogIterative_11_66_0_300_Freq300_uid9
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => logIn_c0,
                 R => lnX_c11);
   FPPow_11_52_Freq300_uid2mult: FPMult_11_66_uid81_Freq300_uid82
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 X => lnX_c11,
                 Y => Y,
                 R => P_c14);
   FPPow_11_52_Freq300_uid2exp: FPExp_11_52_Freq300_uid1477
      port map ( clk  => clk,
                 ce_15 => ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 X => P_c14,
                 R => E_c28);
   flagsE_c28 <= E_c28(wE+wF+2 downto wE+wF+1);
   RisZeroFromExp_c28 <= '1' when flagsE_c28="00" else '0';
   RisZero_c28 <= RisZeroSpecialCase_c28 or RisZeroFromExp_c28;
   RisInfFromExp_c28  <= '1' when flagsE_c28="10" else '0';
   RisInf_c28  <= RisInfSpecialCase_c28 or RisInfFromExp_c28;
   flagR_c28 <= 
           "11" when RisNaN_c28='1'
      else "00" when RisZero_c28='1'
      else "10" when RisInf_c28='1'
      else "01";
   R_expfrac_c28 <= CONV_STD_LOGIC_VECTOR(1023,11) &  CONV_STD_LOGIC_VECTOR(0, 52) when RisOne_c28='1'
       else E_c28(62 downto 0);
   R <= flagR_c28 & signR_c28 & R_expfrac_c28;
end architecture;



