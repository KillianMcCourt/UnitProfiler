--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid17
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid17 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid17 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid22
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid22 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid22 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid27
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid32
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid37
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid37 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid37 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid42
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid42 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid47
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid47 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid47 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid52
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid52 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid52 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid63
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid68
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid73
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid73 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid73 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid78
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid78 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid78 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid83
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid88
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid88 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid88 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid93
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid98
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid113
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid113 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid113 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid118
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid118 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid118 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid123
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid128
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid133
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid133 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid133 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid138
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid143
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid143 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid143 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid148
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid148 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid148 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid153
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid153 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid153 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid158
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid158 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid158 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid163
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid163 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid163 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid168
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid168 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid168 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid183
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid183 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid183 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid188
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid188 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid188 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid193
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid193 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid193 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid198
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid198 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid198 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid203
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid203 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid203 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid208
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid208 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid208 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid213
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid213 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid213 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid218
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid223
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid223 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid223 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid228
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid228 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid228 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid233
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid233 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid233 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid238
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid238 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid238 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid253
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid253 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid253 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid258
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid258 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid258 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid263
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid263 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid263 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid268
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid268 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid268 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid273
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid273 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid273 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid278
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid278 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid278 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid283
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid283 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid283 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid288
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid288 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid288 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid293
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid293 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid293 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid298
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid298 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid298 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid303
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid303 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid303 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid308
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid308 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid308 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid313
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid313 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid313 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid318
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid318 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid318 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq800_uid322
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq800_uid322 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq800_uid322 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq800_uid326
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq800_uid326 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq800_uid326 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq800_uid334
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq800_uid334 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq800_uid334 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq800_uid400
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq800_uid400 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq800_uid400 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq800_uid432
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq800_uid432 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq800_uid432 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid9
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid9 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid9 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid11
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid11 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid11 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid13
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid13 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid13 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid15
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid15 is
   component MultTable_Freq800_uid17 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy18_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid17
      port map ( X => Xtable_c0,
                 Y => Y1_copy18_c0);
   Y1_c0 <= Y1_copy18_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid20
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid20 is
   component MultTable_Freq800_uid22 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy23_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid22
      port map ( X => Xtable_c0,
                 Y => Y1_copy23_c0);
   Y1_c0 <= Y1_copy23_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid25
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid25 is
   component MultTable_Freq800_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid30
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid30 is
   component MultTable_Freq800_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid35
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid35 is
   component MultTable_Freq800_uid37 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy38_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid37
      port map ( X => Xtable_c0,
                 Y => Y1_copy38_c0);
   Y1_c0 <= Y1_copy38_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid40
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid40 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid40 is
   component MultTable_Freq800_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy43_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid42
      port map ( X => Xtable_c0,
                 Y => Y1_copy43_c0);
   Y1_c0 <= Y1_copy43_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid45
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid45 is
   component MultTable_Freq800_uid47 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy48_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid47
      port map ( X => Xtable_c0,
                 Y => Y1_copy48_c0);
   Y1_c0 <= Y1_copy48_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid50
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid50 is
   component MultTable_Freq800_uid52 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy53_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid52
      port map ( X => Xtable_c0,
                 Y => Y1_copy53_c0);
   Y1_c0 <= Y1_copy53_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid55
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid55 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid55 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid57
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid57 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid57 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid59
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid59 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid59 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid61
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid61 is
   component MultTable_Freq800_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid66
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid66 is
   component MultTable_Freq800_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid71
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid71 is
   component MultTable_Freq800_uid73 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy74_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid73
      port map ( X => Xtable_c0,
                 Y => Y1_copy74_c0);
   Y1_c0 <= Y1_copy74_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid76
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid76 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid76 is
   component MultTable_Freq800_uid78 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy79_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid78
      port map ( X => Xtable_c0,
                 Y => Y1_copy79_c0);
   Y1_c0 <= Y1_copy79_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid81
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid81 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid81 is
   component MultTable_Freq800_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy84_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid83
      port map ( X => Xtable_c0,
                 Y => Y1_copy84_c0);
   Y1_c0 <= Y1_copy84_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid86
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid86 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid86 is
   component MultTable_Freq800_uid88 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy89_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid88
      port map ( X => Xtable_c0,
                 Y => Y1_copy89_c0);
   Y1_c0 <= Y1_copy89_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid91
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid91 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid91 is
   component MultTable_Freq800_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid93
      port map ( X => Xtable_c0,
                 Y => Y1_copy94_c0);
   Y1_c0 <= Y1_copy94_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid96
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid96 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid96 is
   component MultTable_Freq800_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid98
      port map ( X => Xtable_c0,
                 Y => Y1_copy99_c0);
   Y1_c0 <= Y1_copy99_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid101
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid101 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid101 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid103
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid103 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid103 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid105
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid105 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid105 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid107
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid107 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid109
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid109 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid111
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid111 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid111 is
   component MultTable_Freq800_uid113 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy114_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid113
      port map ( X => Xtable_c0,
                 Y => Y1_copy114_c0);
   Y1_c0 <= Y1_copy114_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid116
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid116 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid116 is
   component MultTable_Freq800_uid118 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy119_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid118
      port map ( X => Xtable_c0,
                 Y => Y1_copy119_c0);
   Y1_c0 <= Y1_copy119_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid121
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid121 is
   component MultTable_Freq800_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid126
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid126 is
   component MultTable_Freq800_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid131
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid131 is
   component MultTable_Freq800_uid133 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy134_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid133
      port map ( X => Xtable_c0,
                 Y => Y1_copy134_c0);
   Y1_c0 <= Y1_copy134_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid136
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid136 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid136 is
   component MultTable_Freq800_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid138
      port map ( X => Xtable_c0,
                 Y => Y1_copy139_c0);
   Y1_c0 <= Y1_copy139_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid141
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid141 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid141 is
   component MultTable_Freq800_uid143 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy144_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid143
      port map ( X => Xtable_c0,
                 Y => Y1_copy144_c0);
   Y1_c0 <= Y1_copy144_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid146
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid146 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid146 is
   component MultTable_Freq800_uid148 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy149_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid148
      port map ( X => Xtable_c0,
                 Y => Y1_copy149_c0);
   Y1_c0 <= Y1_copy149_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid151
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid151 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid151 is
   component MultTable_Freq800_uid153 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy154_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid153
      port map ( X => Xtable_c0,
                 Y => Y1_copy154_c0);
   Y1_c0 <= Y1_copy154_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid156
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid156 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid156 is
   component MultTable_Freq800_uid158 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy159_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid158
      port map ( X => Xtable_c0,
                 Y => Y1_copy159_c0);
   Y1_c0 <= Y1_copy159_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid161
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid161 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid161 is
   component MultTable_Freq800_uid163 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy164_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid163
      port map ( X => Xtable_c0,
                 Y => Y1_copy164_c0);
   Y1_c0 <= Y1_copy164_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid166
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid166 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid166 is
   component MultTable_Freq800_uid168 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy169_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid168
      port map ( X => Xtable_c0,
                 Y => Y1_copy169_c0);
   Y1_c0 <= Y1_copy169_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid171
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid171 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid171 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid173
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid173 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid173 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid175
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid175 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid175 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid177
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid177 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid177 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid179
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid179 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid179 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid181
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid181 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid181 is
   component MultTable_Freq800_uid183 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy184_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid183
      port map ( X => Xtable_c0,
                 Y => Y1_copy184_c0);
   Y1_c0 <= Y1_copy184_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid186
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid186 is
   component MultTable_Freq800_uid188 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy189_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid188
      port map ( X => Xtable_c0,
                 Y => Y1_copy189_c0);
   Y1_c0 <= Y1_copy189_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid191
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid191 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid191 is
   component MultTable_Freq800_uid193 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy194_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid193
      port map ( X => Xtable_c0,
                 Y => Y1_copy194_c0);
   Y1_c0 <= Y1_copy194_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid196
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid196 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid196 is
   component MultTable_Freq800_uid198 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy199_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid198
      port map ( X => Xtable_c0,
                 Y => Y1_copy199_c0);
   Y1_c0 <= Y1_copy199_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid201
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid201 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid201 is
   component MultTable_Freq800_uid203 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy204_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid203
      port map ( X => Xtable_c0,
                 Y => Y1_copy204_c0);
   Y1_c0 <= Y1_copy204_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid206
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid206 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid206 is
   component MultTable_Freq800_uid208 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy209_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid208
      port map ( X => Xtable_c0,
                 Y => Y1_copy209_c0);
   Y1_c0 <= Y1_copy209_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid211
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid211 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid211 is
   component MultTable_Freq800_uid213 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy214_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid213
      port map ( X => Xtable_c0,
                 Y => Y1_copy214_c0);
   Y1_c0 <= Y1_copy214_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid216
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid216 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid216 is
   component MultTable_Freq800_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid218
      port map ( X => Xtable_c0,
                 Y => Y1_copy219_c0);
   Y1_c0 <= Y1_copy219_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid221
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid221 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid221 is
   component MultTable_Freq800_uid223 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy224_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid223
      port map ( X => Xtable_c0,
                 Y => Y1_copy224_c0);
   Y1_c0 <= Y1_copy224_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid226
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid226 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid226 is
   component MultTable_Freq800_uid228 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy229_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid228
      port map ( X => Xtable_c0,
                 Y => Y1_copy229_c0);
   Y1_c0 <= Y1_copy229_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid231
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid231 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid231 is
   component MultTable_Freq800_uid233 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy234_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid233
      port map ( X => Xtable_c0,
                 Y => Y1_copy234_c0);
   Y1_c0 <= Y1_copy234_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid236
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid236 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid236 is
   component MultTable_Freq800_uid238 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy239_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid238
      port map ( X => Xtable_c0,
                 Y => Y1_copy239_c0);
   Y1_c0 <= Y1_copy239_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid241
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid241 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid241 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid243
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid243 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid243 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid245
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid245 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid245 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid247
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid247 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid247 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid249
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid249 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid249 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid251
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid251 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid251 is
   component MultTable_Freq800_uid253 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy254_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid253
      port map ( X => Xtable_c0,
                 Y => Y1_copy254_c0);
   Y1_c0 <= Y1_copy254_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid256
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid256 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid256 is
   component MultTable_Freq800_uid258 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy259_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid258
      port map ( X => Xtable_c0,
                 Y => Y1_copy259_c0);
   Y1_c0 <= Y1_copy259_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid261
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid261 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid261 is
   component MultTable_Freq800_uid263 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy264_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid263
      port map ( X => Xtable_c0,
                 Y => Y1_copy264_c0);
   Y1_c0 <= Y1_copy264_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid266
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid266 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid266 is
   component MultTable_Freq800_uid268 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy269_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid268
      port map ( X => Xtable_c0,
                 Y => Y1_copy269_c0);
   Y1_c0 <= Y1_copy269_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid271
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid271 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid271 is
   component MultTable_Freq800_uid273 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy274_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid273
      port map ( X => Xtable_c0,
                 Y => Y1_copy274_c0);
   Y1_c0 <= Y1_copy274_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid276
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid276 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid276 is
   component MultTable_Freq800_uid278 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy279_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid278
      port map ( X => Xtable_c0,
                 Y => Y1_copy279_c0);
   Y1_c0 <= Y1_copy279_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid281
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid281 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid281 is
   component MultTable_Freq800_uid283 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy284_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid283
      port map ( X => Xtable_c0,
                 Y => Y1_copy284_c0);
   Y1_c0 <= Y1_copy284_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid286
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid286 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid286 is
   component MultTable_Freq800_uid288 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy289_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid288
      port map ( X => Xtable_c0,
                 Y => Y1_copy289_c0);
   Y1_c0 <= Y1_copy289_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid291
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid291 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid291 is
   component MultTable_Freq800_uid293 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy294_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid293
      port map ( X => Xtable_c0,
                 Y => Y1_copy294_c0);
   Y1_c0 <= Y1_copy294_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid296
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid296 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid296 is
   component MultTable_Freq800_uid298 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy299_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid298
      port map ( X => Xtable_c0,
                 Y => Y1_copy299_c0);
   Y1_c0 <= Y1_copy299_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid301
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid301 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid301 is
   component MultTable_Freq800_uid303 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy304_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid303
      port map ( X => Xtable_c0,
                 Y => Y1_copy304_c0);
   Y1_c0 <= Y1_copy304_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid306
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid306 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid306 is
   component MultTable_Freq800_uid308 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy309_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid308
      port map ( X => Xtable_c0,
                 Y => Y1_copy309_c0);
   Y1_c0 <= Y1_copy309_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid311
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid311 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid311 is
   component MultTable_Freq800_uid313 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy314_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid313
      port map ( X => Xtable_c0,
                 Y => Y1_copy314_c0);
   Y1_c0 <= Y1_copy314_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x3_Freq800_uid316
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid316 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid316 is
   component MultTable_Freq800_uid318 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy319_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid318
      port map ( X => Xtable_c0,
                 Y => Y1_copy319_c0);
   Y1_c0 <= Y1_copy319_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_84_Freq800_uid972
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_84_Freq800_uid972 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
          X : in  std_logic_vector(83 downto 0);
          Y : in  std_logic_vector(83 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(83 downto 0)   );
end entity;

architecture arch of IntAdder_84_Freq800_uid972 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5 :  std_logic;
signal X_0_c4, X_0_c5 :  std_logic_vector(3 downto 0);
signal Y_0_c4, Y_0_c5 :  std_logic_vector(3 downto 0);
signal S_0_c5 :  std_logic_vector(3 downto 0);
signal R_0_c5, R_0_c6, R_0_c7, R_0_c8, R_0_c9, R_0_c10, R_0_c11, R_0_c12, R_0_c13, R_0_c14, R_0_c15, R_0_c16, R_0_c17, R_0_c18, R_0_c19, R_0_c20, R_0_c21, R_0_c22, R_0_c23, R_0_c24, R_0_c25, R_0_c26, R_0_c27, R_0_c28, R_0_c29, R_0_c30, R_0_c31, R_0_c32, R_0_c33 :  std_logic_vector(2 downto 0);
signal Cin_1_c5, Cin_1_c6 :  std_logic;
signal X_1_c4, X_1_c5, X_1_c6 :  std_logic_vector(3 downto 0);
signal Y_1_c4, Y_1_c5, Y_1_c6 :  std_logic_vector(3 downto 0);
signal S_1_c6 :  std_logic_vector(3 downto 0);
signal R_1_c6, R_1_c7, R_1_c8, R_1_c9, R_1_c10, R_1_c11, R_1_c12, R_1_c13, R_1_c14, R_1_c15, R_1_c16, R_1_c17, R_1_c18, R_1_c19, R_1_c20, R_1_c21, R_1_c22, R_1_c23, R_1_c24, R_1_c25, R_1_c26, R_1_c27, R_1_c28, R_1_c29, R_1_c30, R_1_c31, R_1_c32, R_1_c33 :  std_logic_vector(2 downto 0);
signal Cin_2_c6, Cin_2_c7 :  std_logic;
signal X_2_c4, X_2_c5, X_2_c6, X_2_c7 :  std_logic_vector(3 downto 0);
signal Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7 :  std_logic_vector(3 downto 0);
signal S_2_c7 :  std_logic_vector(3 downto 0);
signal R_2_c7, R_2_c8, R_2_c9, R_2_c10, R_2_c11, R_2_c12, R_2_c13, R_2_c14, R_2_c15, R_2_c16, R_2_c17, R_2_c18, R_2_c19, R_2_c20, R_2_c21, R_2_c22, R_2_c23, R_2_c24, R_2_c25, R_2_c26, R_2_c27, R_2_c28, R_2_c29, R_2_c30, R_2_c31, R_2_c32, R_2_c33 :  std_logic_vector(2 downto 0);
signal Cin_3_c7, Cin_3_c8 :  std_logic;
signal X_3_c4, X_3_c5, X_3_c6, X_3_c7, X_3_c8 :  std_logic_vector(3 downto 0);
signal Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8 :  std_logic_vector(3 downto 0);
signal S_3_c8 :  std_logic_vector(3 downto 0);
signal R_3_c8, R_3_c9, R_3_c10, R_3_c11, R_3_c12, R_3_c13, R_3_c14, R_3_c15, R_3_c16, R_3_c17, R_3_c18, R_3_c19, R_3_c20, R_3_c21, R_3_c22, R_3_c23, R_3_c24, R_3_c25, R_3_c26, R_3_c27, R_3_c28, R_3_c29, R_3_c30, R_3_c31, R_3_c32, R_3_c33 :  std_logic_vector(2 downto 0);
signal Cin_4_c8, Cin_4_c9 :  std_logic;
signal X_4_c4, X_4_c5, X_4_c6, X_4_c7, X_4_c8, X_4_c9 :  std_logic_vector(3 downto 0);
signal Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9 :  std_logic_vector(3 downto 0);
signal S_4_c9 :  std_logic_vector(3 downto 0);
signal R_4_c9, R_4_c10, R_4_c11, R_4_c12, R_4_c13, R_4_c14, R_4_c15, R_4_c16, R_4_c17, R_4_c18, R_4_c19, R_4_c20, R_4_c21, R_4_c22, R_4_c23, R_4_c24, R_4_c25, R_4_c26, R_4_c27, R_4_c28, R_4_c29, R_4_c30, R_4_c31, R_4_c32, R_4_c33 :  std_logic_vector(2 downto 0);
signal Cin_5_c9, Cin_5_c10 :  std_logic;
signal X_5_c4, X_5_c5, X_5_c6, X_5_c7, X_5_c8, X_5_c9, X_5_c10 :  std_logic_vector(3 downto 0);
signal Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10 :  std_logic_vector(3 downto 0);
signal S_5_c10 :  std_logic_vector(3 downto 0);
signal R_5_c10, R_5_c11, R_5_c12, R_5_c13, R_5_c14, R_5_c15, R_5_c16, R_5_c17, R_5_c18, R_5_c19, R_5_c20, R_5_c21, R_5_c22, R_5_c23, R_5_c24, R_5_c25, R_5_c26, R_5_c27, R_5_c28, R_5_c29, R_5_c30, R_5_c31, R_5_c32, R_5_c33 :  std_logic_vector(2 downto 0);
signal Cin_6_c10, Cin_6_c11 :  std_logic;
signal X_6_c4, X_6_c5, X_6_c6, X_6_c7, X_6_c8, X_6_c9, X_6_c10, X_6_c11 :  std_logic_vector(3 downto 0);
signal Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11 :  std_logic_vector(3 downto 0);
signal S_6_c11 :  std_logic_vector(3 downto 0);
signal R_6_c11, R_6_c12, R_6_c13, R_6_c14, R_6_c15, R_6_c16, R_6_c17, R_6_c18, R_6_c19, R_6_c20, R_6_c21, R_6_c22, R_6_c23, R_6_c24, R_6_c25, R_6_c26, R_6_c27, R_6_c28, R_6_c29, R_6_c30, R_6_c31, R_6_c32, R_6_c33 :  std_logic_vector(2 downto 0);
signal Cin_7_c11, Cin_7_c12 :  std_logic;
signal X_7_c4, X_7_c5, X_7_c6, X_7_c7, X_7_c8, X_7_c9, X_7_c10, X_7_c11, X_7_c12 :  std_logic_vector(3 downto 0);
signal Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12 :  std_logic_vector(3 downto 0);
signal S_7_c12 :  std_logic_vector(3 downto 0);
signal R_7_c12, R_7_c13, R_7_c14, R_7_c15, R_7_c16, R_7_c17, R_7_c18, R_7_c19, R_7_c20, R_7_c21, R_7_c22, R_7_c23, R_7_c24, R_7_c25, R_7_c26, R_7_c27, R_7_c28, R_7_c29, R_7_c30, R_7_c31, R_7_c32, R_7_c33 :  std_logic_vector(2 downto 0);
signal Cin_8_c12, Cin_8_c13 :  std_logic;
signal X_8_c4, X_8_c5, X_8_c6, X_8_c7, X_8_c8, X_8_c9, X_8_c10, X_8_c11, X_8_c12, X_8_c13 :  std_logic_vector(3 downto 0);
signal Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13 :  std_logic_vector(3 downto 0);
signal S_8_c13 :  std_logic_vector(3 downto 0);
signal R_8_c13, R_8_c14, R_8_c15, R_8_c16, R_8_c17, R_8_c18, R_8_c19, R_8_c20, R_8_c21, R_8_c22, R_8_c23, R_8_c24, R_8_c25, R_8_c26, R_8_c27, R_8_c28, R_8_c29, R_8_c30, R_8_c31, R_8_c32, R_8_c33 :  std_logic_vector(2 downto 0);
signal Cin_9_c13, Cin_9_c14 :  std_logic;
signal X_9_c4, X_9_c5, X_9_c6, X_9_c7, X_9_c8, X_9_c9, X_9_c10, X_9_c11, X_9_c12, X_9_c13, X_9_c14 :  std_logic_vector(3 downto 0);
signal Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14 :  std_logic_vector(3 downto 0);
signal S_9_c14 :  std_logic_vector(3 downto 0);
signal R_9_c14, R_9_c15, R_9_c16, R_9_c17, R_9_c18, R_9_c19, R_9_c20, R_9_c21, R_9_c22, R_9_c23, R_9_c24, R_9_c25, R_9_c26, R_9_c27, R_9_c28, R_9_c29, R_9_c30, R_9_c31, R_9_c32, R_9_c33 :  std_logic_vector(2 downto 0);
signal Cin_10_c14, Cin_10_c15 :  std_logic;
signal X_10_c4, X_10_c5, X_10_c6, X_10_c7, X_10_c8, X_10_c9, X_10_c10, X_10_c11, X_10_c12, X_10_c13, X_10_c14, X_10_c15 :  std_logic_vector(3 downto 0);
signal Y_10_c4, Y_10_c5, Y_10_c6, Y_10_c7, Y_10_c8, Y_10_c9, Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15 :  std_logic_vector(3 downto 0);
signal S_10_c15 :  std_logic_vector(3 downto 0);
signal R_10_c15, R_10_c16, R_10_c17, R_10_c18, R_10_c19, R_10_c20, R_10_c21, R_10_c22, R_10_c23, R_10_c24, R_10_c25, R_10_c26, R_10_c27, R_10_c28, R_10_c29, R_10_c30, R_10_c31, R_10_c32, R_10_c33 :  std_logic_vector(2 downto 0);
signal Cin_11_c15, Cin_11_c16 :  std_logic;
signal X_11_c4, X_11_c5, X_11_c6, X_11_c7, X_11_c8, X_11_c9, X_11_c10, X_11_c11, X_11_c12, X_11_c13, X_11_c14, X_11_c15, X_11_c16 :  std_logic_vector(3 downto 0);
signal Y_11_c4, Y_11_c5, Y_11_c6, Y_11_c7, Y_11_c8, Y_11_c9, Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16 :  std_logic_vector(3 downto 0);
signal S_11_c16 :  std_logic_vector(3 downto 0);
signal R_11_c16, R_11_c17, R_11_c18, R_11_c19, R_11_c20, R_11_c21, R_11_c22, R_11_c23, R_11_c24, R_11_c25, R_11_c26, R_11_c27, R_11_c28, R_11_c29, R_11_c30, R_11_c31, R_11_c32, R_11_c33 :  std_logic_vector(2 downto 0);
signal Cin_12_c16, Cin_12_c17 :  std_logic;
signal X_12_c4, X_12_c5, X_12_c6, X_12_c7, X_12_c8, X_12_c9, X_12_c10, X_12_c11, X_12_c12, X_12_c13, X_12_c14, X_12_c15, X_12_c16, X_12_c17 :  std_logic_vector(3 downto 0);
signal Y_12_c4, Y_12_c5, Y_12_c6, Y_12_c7, Y_12_c8, Y_12_c9, Y_12_c10, Y_12_c11, Y_12_c12, Y_12_c13, Y_12_c14, Y_12_c15, Y_12_c16, Y_12_c17 :  std_logic_vector(3 downto 0);
signal S_12_c17 :  std_logic_vector(3 downto 0);
signal R_12_c17, R_12_c18, R_12_c19, R_12_c20, R_12_c21, R_12_c22, R_12_c23, R_12_c24, R_12_c25, R_12_c26, R_12_c27, R_12_c28, R_12_c29, R_12_c30, R_12_c31, R_12_c32, R_12_c33 :  std_logic_vector(2 downto 0);
signal Cin_13_c17, Cin_13_c18 :  std_logic;
signal X_13_c4, X_13_c5, X_13_c6, X_13_c7, X_13_c8, X_13_c9, X_13_c10, X_13_c11, X_13_c12, X_13_c13, X_13_c14, X_13_c15, X_13_c16, X_13_c17, X_13_c18 :  std_logic_vector(3 downto 0);
signal Y_13_c4, Y_13_c5, Y_13_c6, Y_13_c7, Y_13_c8, Y_13_c9, Y_13_c10, Y_13_c11, Y_13_c12, Y_13_c13, Y_13_c14, Y_13_c15, Y_13_c16, Y_13_c17, Y_13_c18 :  std_logic_vector(3 downto 0);
signal S_13_c18 :  std_logic_vector(3 downto 0);
signal R_13_c18, R_13_c19, R_13_c20, R_13_c21, R_13_c22, R_13_c23, R_13_c24, R_13_c25, R_13_c26, R_13_c27, R_13_c28, R_13_c29, R_13_c30, R_13_c31, R_13_c32, R_13_c33 :  std_logic_vector(2 downto 0);
signal Cin_14_c18, Cin_14_c19, Cin_14_c20 :  std_logic;
signal X_14_c4, X_14_c5, X_14_c6, X_14_c7, X_14_c8, X_14_c9, X_14_c10, X_14_c11, X_14_c12, X_14_c13, X_14_c14, X_14_c15, X_14_c16, X_14_c17, X_14_c18, X_14_c19, X_14_c20 :  std_logic_vector(3 downto 0);
signal Y_14_c4, Y_14_c5, Y_14_c6, Y_14_c7, Y_14_c8, Y_14_c9, Y_14_c10, Y_14_c11, Y_14_c12, Y_14_c13, Y_14_c14, Y_14_c15, Y_14_c16, Y_14_c17, Y_14_c18, Y_14_c19, Y_14_c20 :  std_logic_vector(3 downto 0);
signal S_14_c20 :  std_logic_vector(3 downto 0);
signal R_14_c20, R_14_c21, R_14_c22, R_14_c23, R_14_c24, R_14_c25, R_14_c26, R_14_c27, R_14_c28, R_14_c29, R_14_c30, R_14_c31, R_14_c32, R_14_c33 :  std_logic_vector(2 downto 0);
signal Cin_15_c20, Cin_15_c21 :  std_logic;
signal X_15_c4, X_15_c5, X_15_c6, X_15_c7, X_15_c8, X_15_c9, X_15_c10, X_15_c11, X_15_c12, X_15_c13, X_15_c14, X_15_c15, X_15_c16, X_15_c17, X_15_c18, X_15_c19, X_15_c20, X_15_c21 :  std_logic_vector(3 downto 0);
signal Y_15_c4, Y_15_c5, Y_15_c6, Y_15_c7, Y_15_c8, Y_15_c9, Y_15_c10, Y_15_c11, Y_15_c12, Y_15_c13, Y_15_c14, Y_15_c15, Y_15_c16, Y_15_c17, Y_15_c18, Y_15_c19, Y_15_c20, Y_15_c21 :  std_logic_vector(3 downto 0);
signal S_15_c21 :  std_logic_vector(3 downto 0);
signal R_15_c21, R_15_c22, R_15_c23, R_15_c24, R_15_c25, R_15_c26, R_15_c27, R_15_c28, R_15_c29, R_15_c30, R_15_c31, R_15_c32, R_15_c33 :  std_logic_vector(2 downto 0);
signal Cin_16_c21, Cin_16_c22 :  std_logic;
signal X_16_c4, X_16_c5, X_16_c6, X_16_c7, X_16_c8, X_16_c9, X_16_c10, X_16_c11, X_16_c12, X_16_c13, X_16_c14, X_16_c15, X_16_c16, X_16_c17, X_16_c18, X_16_c19, X_16_c20, X_16_c21, X_16_c22 :  std_logic_vector(3 downto 0);
signal Y_16_c4, Y_16_c5, Y_16_c6, Y_16_c7, Y_16_c8, Y_16_c9, Y_16_c10, Y_16_c11, Y_16_c12, Y_16_c13, Y_16_c14, Y_16_c15, Y_16_c16, Y_16_c17, Y_16_c18, Y_16_c19, Y_16_c20, Y_16_c21, Y_16_c22 :  std_logic_vector(3 downto 0);
signal S_16_c22 :  std_logic_vector(3 downto 0);
signal R_16_c22, R_16_c23, R_16_c24, R_16_c25, R_16_c26, R_16_c27, R_16_c28, R_16_c29, R_16_c30, R_16_c31, R_16_c32, R_16_c33 :  std_logic_vector(2 downto 0);
signal Cin_17_c22, Cin_17_c23 :  std_logic;
signal X_17_c4, X_17_c5, X_17_c6, X_17_c7, X_17_c8, X_17_c9, X_17_c10, X_17_c11, X_17_c12, X_17_c13, X_17_c14, X_17_c15, X_17_c16, X_17_c17, X_17_c18, X_17_c19, X_17_c20, X_17_c21, X_17_c22, X_17_c23 :  std_logic_vector(3 downto 0);
signal Y_17_c4, Y_17_c5, Y_17_c6, Y_17_c7, Y_17_c8, Y_17_c9, Y_17_c10, Y_17_c11, Y_17_c12, Y_17_c13, Y_17_c14, Y_17_c15, Y_17_c16, Y_17_c17, Y_17_c18, Y_17_c19, Y_17_c20, Y_17_c21, Y_17_c22, Y_17_c23 :  std_logic_vector(3 downto 0);
signal S_17_c23 :  std_logic_vector(3 downto 0);
signal R_17_c23, R_17_c24, R_17_c25, R_17_c26, R_17_c27, R_17_c28, R_17_c29, R_17_c30, R_17_c31, R_17_c32, R_17_c33 :  std_logic_vector(2 downto 0);
signal Cin_18_c23, Cin_18_c24 :  std_logic;
signal X_18_c4, X_18_c5, X_18_c6, X_18_c7, X_18_c8, X_18_c9, X_18_c10, X_18_c11, X_18_c12, X_18_c13, X_18_c14, X_18_c15, X_18_c16, X_18_c17, X_18_c18, X_18_c19, X_18_c20, X_18_c21, X_18_c22, X_18_c23, X_18_c24 :  std_logic_vector(3 downto 0);
signal Y_18_c4, Y_18_c5, Y_18_c6, Y_18_c7, Y_18_c8, Y_18_c9, Y_18_c10, Y_18_c11, Y_18_c12, Y_18_c13, Y_18_c14, Y_18_c15, Y_18_c16, Y_18_c17, Y_18_c18, Y_18_c19, Y_18_c20, Y_18_c21, Y_18_c22, Y_18_c23, Y_18_c24 :  std_logic_vector(3 downto 0);
signal S_18_c24 :  std_logic_vector(3 downto 0);
signal R_18_c24, R_18_c25, R_18_c26, R_18_c27, R_18_c28, R_18_c29, R_18_c30, R_18_c31, R_18_c32, R_18_c33 :  std_logic_vector(2 downto 0);
signal Cin_19_c24, Cin_19_c25 :  std_logic;
signal X_19_c4, X_19_c5, X_19_c6, X_19_c7, X_19_c8, X_19_c9, X_19_c10, X_19_c11, X_19_c12, X_19_c13, X_19_c14, X_19_c15, X_19_c16, X_19_c17, X_19_c18, X_19_c19, X_19_c20, X_19_c21, X_19_c22, X_19_c23, X_19_c24, X_19_c25 :  std_logic_vector(3 downto 0);
signal Y_19_c4, Y_19_c5, Y_19_c6, Y_19_c7, Y_19_c8, Y_19_c9, Y_19_c10, Y_19_c11, Y_19_c12, Y_19_c13, Y_19_c14, Y_19_c15, Y_19_c16, Y_19_c17, Y_19_c18, Y_19_c19, Y_19_c20, Y_19_c21, Y_19_c22, Y_19_c23, Y_19_c24, Y_19_c25 :  std_logic_vector(3 downto 0);
signal S_19_c25 :  std_logic_vector(3 downto 0);
signal R_19_c25, R_19_c26, R_19_c27, R_19_c28, R_19_c29, R_19_c30, R_19_c31, R_19_c32, R_19_c33 :  std_logic_vector(2 downto 0);
signal Cin_20_c25, Cin_20_c26 :  std_logic;
signal X_20_c4, X_20_c5, X_20_c6, X_20_c7, X_20_c8, X_20_c9, X_20_c10, X_20_c11, X_20_c12, X_20_c13, X_20_c14, X_20_c15, X_20_c16, X_20_c17, X_20_c18, X_20_c19, X_20_c20, X_20_c21, X_20_c22, X_20_c23, X_20_c24, X_20_c25, X_20_c26 :  std_logic_vector(3 downto 0);
signal Y_20_c4, Y_20_c5, Y_20_c6, Y_20_c7, Y_20_c8, Y_20_c9, Y_20_c10, Y_20_c11, Y_20_c12, Y_20_c13, Y_20_c14, Y_20_c15, Y_20_c16, Y_20_c17, Y_20_c18, Y_20_c19, Y_20_c20, Y_20_c21, Y_20_c22, Y_20_c23, Y_20_c24, Y_20_c25, Y_20_c26 :  std_logic_vector(3 downto 0);
signal S_20_c26 :  std_logic_vector(3 downto 0);
signal R_20_c26, R_20_c27, R_20_c28, R_20_c29, R_20_c30, R_20_c31, R_20_c32, R_20_c33 :  std_logic_vector(2 downto 0);
signal Cin_21_c26, Cin_21_c27 :  std_logic;
signal X_21_c4, X_21_c5, X_21_c6, X_21_c7, X_21_c8, X_21_c9, X_21_c10, X_21_c11, X_21_c12, X_21_c13, X_21_c14, X_21_c15, X_21_c16, X_21_c17, X_21_c18, X_21_c19, X_21_c20, X_21_c21, X_21_c22, X_21_c23, X_21_c24, X_21_c25, X_21_c26, X_21_c27 :  std_logic_vector(3 downto 0);
signal Y_21_c4, Y_21_c5, Y_21_c6, Y_21_c7, Y_21_c8, Y_21_c9, Y_21_c10, Y_21_c11, Y_21_c12, Y_21_c13, Y_21_c14, Y_21_c15, Y_21_c16, Y_21_c17, Y_21_c18, Y_21_c19, Y_21_c20, Y_21_c21, Y_21_c22, Y_21_c23, Y_21_c24, Y_21_c25, Y_21_c26, Y_21_c27 :  std_logic_vector(3 downto 0);
signal S_21_c27 :  std_logic_vector(3 downto 0);
signal R_21_c27, R_21_c28, R_21_c29, R_21_c30, R_21_c31, R_21_c32, R_21_c33 :  std_logic_vector(2 downto 0);
signal Cin_22_c27, Cin_22_c28 :  std_logic;
signal X_22_c4, X_22_c5, X_22_c6, X_22_c7, X_22_c8, X_22_c9, X_22_c10, X_22_c11, X_22_c12, X_22_c13, X_22_c14, X_22_c15, X_22_c16, X_22_c17, X_22_c18, X_22_c19, X_22_c20, X_22_c21, X_22_c22, X_22_c23, X_22_c24, X_22_c25, X_22_c26, X_22_c27, X_22_c28 :  std_logic_vector(3 downto 0);
signal Y_22_c4, Y_22_c5, Y_22_c6, Y_22_c7, Y_22_c8, Y_22_c9, Y_22_c10, Y_22_c11, Y_22_c12, Y_22_c13, Y_22_c14, Y_22_c15, Y_22_c16, Y_22_c17, Y_22_c18, Y_22_c19, Y_22_c20, Y_22_c21, Y_22_c22, Y_22_c23, Y_22_c24, Y_22_c25, Y_22_c26, Y_22_c27, Y_22_c28 :  std_logic_vector(3 downto 0);
signal S_22_c28 :  std_logic_vector(3 downto 0);
signal R_22_c28, R_22_c29, R_22_c30, R_22_c31, R_22_c32, R_22_c33 :  std_logic_vector(2 downto 0);
signal Cin_23_c28, Cin_23_c29 :  std_logic;
signal X_23_c4, X_23_c5, X_23_c6, X_23_c7, X_23_c8, X_23_c9, X_23_c10, X_23_c11, X_23_c12, X_23_c13, X_23_c14, X_23_c15, X_23_c16, X_23_c17, X_23_c18, X_23_c19, X_23_c20, X_23_c21, X_23_c22, X_23_c23, X_23_c24, X_23_c25, X_23_c26, X_23_c27, X_23_c28, X_23_c29 :  std_logic_vector(3 downto 0);
signal Y_23_c4, Y_23_c5, Y_23_c6, Y_23_c7, Y_23_c8, Y_23_c9, Y_23_c10, Y_23_c11, Y_23_c12, Y_23_c13, Y_23_c14, Y_23_c15, Y_23_c16, Y_23_c17, Y_23_c18, Y_23_c19, Y_23_c20, Y_23_c21, Y_23_c22, Y_23_c23, Y_23_c24, Y_23_c25, Y_23_c26, Y_23_c27, Y_23_c28, Y_23_c29 :  std_logic_vector(3 downto 0);
signal S_23_c29 :  std_logic_vector(3 downto 0);
signal R_23_c29, R_23_c30, R_23_c31, R_23_c32, R_23_c33 :  std_logic_vector(2 downto 0);
signal Cin_24_c29, Cin_24_c30 :  std_logic;
signal X_24_c4, X_24_c5, X_24_c6, X_24_c7, X_24_c8, X_24_c9, X_24_c10, X_24_c11, X_24_c12, X_24_c13, X_24_c14, X_24_c15, X_24_c16, X_24_c17, X_24_c18, X_24_c19, X_24_c20, X_24_c21, X_24_c22, X_24_c23, X_24_c24, X_24_c25, X_24_c26, X_24_c27, X_24_c28, X_24_c29, X_24_c30 :  std_logic_vector(3 downto 0);
signal Y_24_c4, Y_24_c5, Y_24_c6, Y_24_c7, Y_24_c8, Y_24_c9, Y_24_c10, Y_24_c11, Y_24_c12, Y_24_c13, Y_24_c14, Y_24_c15, Y_24_c16, Y_24_c17, Y_24_c18, Y_24_c19, Y_24_c20, Y_24_c21, Y_24_c22, Y_24_c23, Y_24_c24, Y_24_c25, Y_24_c26, Y_24_c27, Y_24_c28, Y_24_c29, Y_24_c30 :  std_logic_vector(3 downto 0);
signal S_24_c30 :  std_logic_vector(3 downto 0);
signal R_24_c30, R_24_c31, R_24_c32, R_24_c33 :  std_logic_vector(2 downto 0);
signal Cin_25_c30, Cin_25_c31 :  std_logic;
signal X_25_c4, X_25_c5, X_25_c6, X_25_c7, X_25_c8, X_25_c9, X_25_c10, X_25_c11, X_25_c12, X_25_c13, X_25_c14, X_25_c15, X_25_c16, X_25_c17, X_25_c18, X_25_c19, X_25_c20, X_25_c21, X_25_c22, X_25_c23, X_25_c24, X_25_c25, X_25_c26, X_25_c27, X_25_c28, X_25_c29, X_25_c30, X_25_c31 :  std_logic_vector(3 downto 0);
signal Y_25_c4, Y_25_c5, Y_25_c6, Y_25_c7, Y_25_c8, Y_25_c9, Y_25_c10, Y_25_c11, Y_25_c12, Y_25_c13, Y_25_c14, Y_25_c15, Y_25_c16, Y_25_c17, Y_25_c18, Y_25_c19, Y_25_c20, Y_25_c21, Y_25_c22, Y_25_c23, Y_25_c24, Y_25_c25, Y_25_c26, Y_25_c27, Y_25_c28, Y_25_c29, Y_25_c30, Y_25_c31 :  std_logic_vector(3 downto 0);
signal S_25_c31 :  std_logic_vector(3 downto 0);
signal R_25_c31, R_25_c32, R_25_c33 :  std_logic_vector(2 downto 0);
signal Cin_26_c31, Cin_26_c32 :  std_logic;
signal X_26_c4, X_26_c5, X_26_c6, X_26_c7, X_26_c8, X_26_c9, X_26_c10, X_26_c11, X_26_c12, X_26_c13, X_26_c14, X_26_c15, X_26_c16, X_26_c17, X_26_c18, X_26_c19, X_26_c20, X_26_c21, X_26_c22, X_26_c23, X_26_c24, X_26_c25, X_26_c26, X_26_c27, X_26_c28, X_26_c29, X_26_c30, X_26_c31, X_26_c32 :  std_logic_vector(3 downto 0);
signal Y_26_c4, Y_26_c5, Y_26_c6, Y_26_c7, Y_26_c8, Y_26_c9, Y_26_c10, Y_26_c11, Y_26_c12, Y_26_c13, Y_26_c14, Y_26_c15, Y_26_c16, Y_26_c17, Y_26_c18, Y_26_c19, Y_26_c20, Y_26_c21, Y_26_c22, Y_26_c23, Y_26_c24, Y_26_c25, Y_26_c26, Y_26_c27, Y_26_c28, Y_26_c29, Y_26_c30, Y_26_c31, Y_26_c32 :  std_logic_vector(3 downto 0);
signal S_26_c32 :  std_logic_vector(3 downto 0);
signal R_26_c32, R_26_c33 :  std_logic_vector(2 downto 0);
signal Cin_27_c32, Cin_27_c33 :  std_logic;
signal X_27_c4, X_27_c5, X_27_c6, X_27_c7, X_27_c8, X_27_c9, X_27_c10, X_27_c11, X_27_c12, X_27_c13, X_27_c14, X_27_c15, X_27_c16, X_27_c17, X_27_c18, X_27_c19, X_27_c20, X_27_c21, X_27_c22, X_27_c23, X_27_c24, X_27_c25, X_27_c26, X_27_c27, X_27_c28, X_27_c29, X_27_c30, X_27_c31, X_27_c32, X_27_c33 :  std_logic_vector(3 downto 0);
signal Y_27_c4, Y_27_c5, Y_27_c6, Y_27_c7, Y_27_c8, Y_27_c9, Y_27_c10, Y_27_c11, Y_27_c12, Y_27_c13, Y_27_c14, Y_27_c15, Y_27_c16, Y_27_c17, Y_27_c18, Y_27_c19, Y_27_c20, Y_27_c21, Y_27_c22, Y_27_c23, Y_27_c24, Y_27_c25, Y_27_c26, Y_27_c27, Y_27_c28, Y_27_c29, Y_27_c30, Y_27_c31, Y_27_c32, Y_27_c33 :  std_logic_vector(3 downto 0);
signal S_27_c33 :  std_logic_vector(3 downto 0);
signal R_27_c33 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
               X_0_c5 <= X_0_c4;
               Y_0_c5 <= Y_0_c4;
               X_1_c5 <= X_1_c4;
               Y_1_c5 <= Y_1_c4;
               X_2_c5 <= X_2_c4;
               Y_2_c5 <= Y_2_c4;
               X_3_c5 <= X_3_c4;
               Y_3_c5 <= Y_3_c4;
               X_4_c5 <= X_4_c4;
               Y_4_c5 <= Y_4_c4;
               X_5_c5 <= X_5_c4;
               Y_5_c5 <= Y_5_c4;
               X_6_c5 <= X_6_c4;
               Y_6_c5 <= Y_6_c4;
               X_7_c5 <= X_7_c4;
               Y_7_c5 <= Y_7_c4;
               X_8_c5 <= X_8_c4;
               Y_8_c5 <= Y_8_c4;
               X_9_c5 <= X_9_c4;
               Y_9_c5 <= Y_9_c4;
               X_10_c5 <= X_10_c4;
               Y_10_c5 <= Y_10_c4;
               X_11_c5 <= X_11_c4;
               Y_11_c5 <= Y_11_c4;
               X_12_c5 <= X_12_c4;
               Y_12_c5 <= Y_12_c4;
               X_13_c5 <= X_13_c4;
               Y_13_c5 <= Y_13_c4;
               X_14_c5 <= X_14_c4;
               Y_14_c5 <= Y_14_c4;
               X_15_c5 <= X_15_c4;
               Y_15_c5 <= Y_15_c4;
               X_16_c5 <= X_16_c4;
               Y_16_c5 <= Y_16_c4;
               X_17_c5 <= X_17_c4;
               Y_17_c5 <= Y_17_c4;
               X_18_c5 <= X_18_c4;
               Y_18_c5 <= Y_18_c4;
               X_19_c5 <= X_19_c4;
               Y_19_c5 <= Y_19_c4;
               X_20_c5 <= X_20_c4;
               Y_20_c5 <= Y_20_c4;
               X_21_c5 <= X_21_c4;
               Y_21_c5 <= Y_21_c4;
               X_22_c5 <= X_22_c4;
               Y_22_c5 <= Y_22_c4;
               X_23_c5 <= X_23_c4;
               Y_23_c5 <= Y_23_c4;
               X_24_c5 <= X_24_c4;
               Y_24_c5 <= Y_24_c4;
               X_25_c5 <= X_25_c4;
               Y_25_c5 <= Y_25_c4;
               X_26_c5 <= X_26_c4;
               Y_26_c5 <= Y_26_c4;
               X_27_c5 <= X_27_c4;
               Y_27_c5 <= Y_27_c4;
            end if;
            if ce_6 = '1' then
               R_0_c6 <= R_0_c5;
               Cin_1_c6 <= Cin_1_c5;
               X_1_c6 <= X_1_c5;
               Y_1_c6 <= Y_1_c5;
               X_2_c6 <= X_2_c5;
               Y_2_c6 <= Y_2_c5;
               X_3_c6 <= X_3_c5;
               Y_3_c6 <= Y_3_c5;
               X_4_c6 <= X_4_c5;
               Y_4_c6 <= Y_4_c5;
               X_5_c6 <= X_5_c5;
               Y_5_c6 <= Y_5_c5;
               X_6_c6 <= X_6_c5;
               Y_6_c6 <= Y_6_c5;
               X_7_c6 <= X_7_c5;
               Y_7_c6 <= Y_7_c5;
               X_8_c6 <= X_8_c5;
               Y_8_c6 <= Y_8_c5;
               X_9_c6 <= X_9_c5;
               Y_9_c6 <= Y_9_c5;
               X_10_c6 <= X_10_c5;
               Y_10_c6 <= Y_10_c5;
               X_11_c6 <= X_11_c5;
               Y_11_c6 <= Y_11_c5;
               X_12_c6 <= X_12_c5;
               Y_12_c6 <= Y_12_c5;
               X_13_c6 <= X_13_c5;
               Y_13_c6 <= Y_13_c5;
               X_14_c6 <= X_14_c5;
               Y_14_c6 <= Y_14_c5;
               X_15_c6 <= X_15_c5;
               Y_15_c6 <= Y_15_c5;
               X_16_c6 <= X_16_c5;
               Y_16_c6 <= Y_16_c5;
               X_17_c6 <= X_17_c5;
               Y_17_c6 <= Y_17_c5;
               X_18_c6 <= X_18_c5;
               Y_18_c6 <= Y_18_c5;
               X_19_c6 <= X_19_c5;
               Y_19_c6 <= Y_19_c5;
               X_20_c6 <= X_20_c5;
               Y_20_c6 <= Y_20_c5;
               X_21_c6 <= X_21_c5;
               Y_21_c6 <= Y_21_c5;
               X_22_c6 <= X_22_c5;
               Y_22_c6 <= Y_22_c5;
               X_23_c6 <= X_23_c5;
               Y_23_c6 <= Y_23_c5;
               X_24_c6 <= X_24_c5;
               Y_24_c6 <= Y_24_c5;
               X_25_c6 <= X_25_c5;
               Y_25_c6 <= Y_25_c5;
               X_26_c6 <= X_26_c5;
               Y_26_c6 <= Y_26_c5;
               X_27_c6 <= X_27_c5;
               Y_27_c6 <= Y_27_c5;
            end if;
            if ce_7 = '1' then
               R_0_c7 <= R_0_c6;
               R_1_c7 <= R_1_c6;
               Cin_2_c7 <= Cin_2_c6;
               X_2_c7 <= X_2_c6;
               Y_2_c7 <= Y_2_c6;
               X_3_c7 <= X_3_c6;
               Y_3_c7 <= Y_3_c6;
               X_4_c7 <= X_4_c6;
               Y_4_c7 <= Y_4_c6;
               X_5_c7 <= X_5_c6;
               Y_5_c7 <= Y_5_c6;
               X_6_c7 <= X_6_c6;
               Y_6_c7 <= Y_6_c6;
               X_7_c7 <= X_7_c6;
               Y_7_c7 <= Y_7_c6;
               X_8_c7 <= X_8_c6;
               Y_8_c7 <= Y_8_c6;
               X_9_c7 <= X_9_c6;
               Y_9_c7 <= Y_9_c6;
               X_10_c7 <= X_10_c6;
               Y_10_c7 <= Y_10_c6;
               X_11_c7 <= X_11_c6;
               Y_11_c7 <= Y_11_c6;
               X_12_c7 <= X_12_c6;
               Y_12_c7 <= Y_12_c6;
               X_13_c7 <= X_13_c6;
               Y_13_c7 <= Y_13_c6;
               X_14_c7 <= X_14_c6;
               Y_14_c7 <= Y_14_c6;
               X_15_c7 <= X_15_c6;
               Y_15_c7 <= Y_15_c6;
               X_16_c7 <= X_16_c6;
               Y_16_c7 <= Y_16_c6;
               X_17_c7 <= X_17_c6;
               Y_17_c7 <= Y_17_c6;
               X_18_c7 <= X_18_c6;
               Y_18_c7 <= Y_18_c6;
               X_19_c7 <= X_19_c6;
               Y_19_c7 <= Y_19_c6;
               X_20_c7 <= X_20_c6;
               Y_20_c7 <= Y_20_c6;
               X_21_c7 <= X_21_c6;
               Y_21_c7 <= Y_21_c6;
               X_22_c7 <= X_22_c6;
               Y_22_c7 <= Y_22_c6;
               X_23_c7 <= X_23_c6;
               Y_23_c7 <= Y_23_c6;
               X_24_c7 <= X_24_c6;
               Y_24_c7 <= Y_24_c6;
               X_25_c7 <= X_25_c6;
               Y_25_c7 <= Y_25_c6;
               X_26_c7 <= X_26_c6;
               Y_26_c7 <= Y_26_c6;
               X_27_c7 <= X_27_c6;
               Y_27_c7 <= Y_27_c6;
            end if;
            if ce_8 = '1' then
               R_0_c8 <= R_0_c7;
               R_1_c8 <= R_1_c7;
               R_2_c8 <= R_2_c7;
               Cin_3_c8 <= Cin_3_c7;
               X_3_c8 <= X_3_c7;
               Y_3_c8 <= Y_3_c7;
               X_4_c8 <= X_4_c7;
               Y_4_c8 <= Y_4_c7;
               X_5_c8 <= X_5_c7;
               Y_5_c8 <= Y_5_c7;
               X_6_c8 <= X_6_c7;
               Y_6_c8 <= Y_6_c7;
               X_7_c8 <= X_7_c7;
               Y_7_c8 <= Y_7_c7;
               X_8_c8 <= X_8_c7;
               Y_8_c8 <= Y_8_c7;
               X_9_c8 <= X_9_c7;
               Y_9_c8 <= Y_9_c7;
               X_10_c8 <= X_10_c7;
               Y_10_c8 <= Y_10_c7;
               X_11_c8 <= X_11_c7;
               Y_11_c8 <= Y_11_c7;
               X_12_c8 <= X_12_c7;
               Y_12_c8 <= Y_12_c7;
               X_13_c8 <= X_13_c7;
               Y_13_c8 <= Y_13_c7;
               X_14_c8 <= X_14_c7;
               Y_14_c8 <= Y_14_c7;
               X_15_c8 <= X_15_c7;
               Y_15_c8 <= Y_15_c7;
               X_16_c8 <= X_16_c7;
               Y_16_c8 <= Y_16_c7;
               X_17_c8 <= X_17_c7;
               Y_17_c8 <= Y_17_c7;
               X_18_c8 <= X_18_c7;
               Y_18_c8 <= Y_18_c7;
               X_19_c8 <= X_19_c7;
               Y_19_c8 <= Y_19_c7;
               X_20_c8 <= X_20_c7;
               Y_20_c8 <= Y_20_c7;
               X_21_c8 <= X_21_c7;
               Y_21_c8 <= Y_21_c7;
               X_22_c8 <= X_22_c7;
               Y_22_c8 <= Y_22_c7;
               X_23_c8 <= X_23_c7;
               Y_23_c8 <= Y_23_c7;
               X_24_c8 <= X_24_c7;
               Y_24_c8 <= Y_24_c7;
               X_25_c8 <= X_25_c7;
               Y_25_c8 <= Y_25_c7;
               X_26_c8 <= X_26_c7;
               Y_26_c8 <= Y_26_c7;
               X_27_c8 <= X_27_c7;
               Y_27_c8 <= Y_27_c7;
            end if;
            if ce_9 = '1' then
               R_0_c9 <= R_0_c8;
               R_1_c9 <= R_1_c8;
               R_2_c9 <= R_2_c8;
               R_3_c9 <= R_3_c8;
               Cin_4_c9 <= Cin_4_c8;
               X_4_c9 <= X_4_c8;
               Y_4_c9 <= Y_4_c8;
               X_5_c9 <= X_5_c8;
               Y_5_c9 <= Y_5_c8;
               X_6_c9 <= X_6_c8;
               Y_6_c9 <= Y_6_c8;
               X_7_c9 <= X_7_c8;
               Y_7_c9 <= Y_7_c8;
               X_8_c9 <= X_8_c8;
               Y_8_c9 <= Y_8_c8;
               X_9_c9 <= X_9_c8;
               Y_9_c9 <= Y_9_c8;
               X_10_c9 <= X_10_c8;
               Y_10_c9 <= Y_10_c8;
               X_11_c9 <= X_11_c8;
               Y_11_c9 <= Y_11_c8;
               X_12_c9 <= X_12_c8;
               Y_12_c9 <= Y_12_c8;
               X_13_c9 <= X_13_c8;
               Y_13_c9 <= Y_13_c8;
               X_14_c9 <= X_14_c8;
               Y_14_c9 <= Y_14_c8;
               X_15_c9 <= X_15_c8;
               Y_15_c9 <= Y_15_c8;
               X_16_c9 <= X_16_c8;
               Y_16_c9 <= Y_16_c8;
               X_17_c9 <= X_17_c8;
               Y_17_c9 <= Y_17_c8;
               X_18_c9 <= X_18_c8;
               Y_18_c9 <= Y_18_c8;
               X_19_c9 <= X_19_c8;
               Y_19_c9 <= Y_19_c8;
               X_20_c9 <= X_20_c8;
               Y_20_c9 <= Y_20_c8;
               X_21_c9 <= X_21_c8;
               Y_21_c9 <= Y_21_c8;
               X_22_c9 <= X_22_c8;
               Y_22_c9 <= Y_22_c8;
               X_23_c9 <= X_23_c8;
               Y_23_c9 <= Y_23_c8;
               X_24_c9 <= X_24_c8;
               Y_24_c9 <= Y_24_c8;
               X_25_c9 <= X_25_c8;
               Y_25_c9 <= Y_25_c8;
               X_26_c9 <= X_26_c8;
               Y_26_c9 <= Y_26_c8;
               X_27_c9 <= X_27_c8;
               Y_27_c9 <= Y_27_c8;
            end if;
            if ce_10 = '1' then
               R_0_c10 <= R_0_c9;
               R_1_c10 <= R_1_c9;
               R_2_c10 <= R_2_c9;
               R_3_c10 <= R_3_c9;
               R_4_c10 <= R_4_c9;
               Cin_5_c10 <= Cin_5_c9;
               X_5_c10 <= X_5_c9;
               Y_5_c10 <= Y_5_c9;
               X_6_c10 <= X_6_c9;
               Y_6_c10 <= Y_6_c9;
               X_7_c10 <= X_7_c9;
               Y_7_c10 <= Y_7_c9;
               X_8_c10 <= X_8_c9;
               Y_8_c10 <= Y_8_c9;
               X_9_c10 <= X_9_c9;
               Y_9_c10 <= Y_9_c9;
               X_10_c10 <= X_10_c9;
               Y_10_c10 <= Y_10_c9;
               X_11_c10 <= X_11_c9;
               Y_11_c10 <= Y_11_c9;
               X_12_c10 <= X_12_c9;
               Y_12_c10 <= Y_12_c9;
               X_13_c10 <= X_13_c9;
               Y_13_c10 <= Y_13_c9;
               X_14_c10 <= X_14_c9;
               Y_14_c10 <= Y_14_c9;
               X_15_c10 <= X_15_c9;
               Y_15_c10 <= Y_15_c9;
               X_16_c10 <= X_16_c9;
               Y_16_c10 <= Y_16_c9;
               X_17_c10 <= X_17_c9;
               Y_17_c10 <= Y_17_c9;
               X_18_c10 <= X_18_c9;
               Y_18_c10 <= Y_18_c9;
               X_19_c10 <= X_19_c9;
               Y_19_c10 <= Y_19_c9;
               X_20_c10 <= X_20_c9;
               Y_20_c10 <= Y_20_c9;
               X_21_c10 <= X_21_c9;
               Y_21_c10 <= Y_21_c9;
               X_22_c10 <= X_22_c9;
               Y_22_c10 <= Y_22_c9;
               X_23_c10 <= X_23_c9;
               Y_23_c10 <= Y_23_c9;
               X_24_c10 <= X_24_c9;
               Y_24_c10 <= Y_24_c9;
               X_25_c10 <= X_25_c9;
               Y_25_c10 <= Y_25_c9;
               X_26_c10 <= X_26_c9;
               Y_26_c10 <= Y_26_c9;
               X_27_c10 <= X_27_c9;
               Y_27_c10 <= Y_27_c9;
            end if;
            if ce_11 = '1' then
               R_0_c11 <= R_0_c10;
               R_1_c11 <= R_1_c10;
               R_2_c11 <= R_2_c10;
               R_3_c11 <= R_3_c10;
               R_4_c11 <= R_4_c10;
               R_5_c11 <= R_5_c10;
               Cin_6_c11 <= Cin_6_c10;
               X_6_c11 <= X_6_c10;
               Y_6_c11 <= Y_6_c10;
               X_7_c11 <= X_7_c10;
               Y_7_c11 <= Y_7_c10;
               X_8_c11 <= X_8_c10;
               Y_8_c11 <= Y_8_c10;
               X_9_c11 <= X_9_c10;
               Y_9_c11 <= Y_9_c10;
               X_10_c11 <= X_10_c10;
               Y_10_c11 <= Y_10_c10;
               X_11_c11 <= X_11_c10;
               Y_11_c11 <= Y_11_c10;
               X_12_c11 <= X_12_c10;
               Y_12_c11 <= Y_12_c10;
               X_13_c11 <= X_13_c10;
               Y_13_c11 <= Y_13_c10;
               X_14_c11 <= X_14_c10;
               Y_14_c11 <= Y_14_c10;
               X_15_c11 <= X_15_c10;
               Y_15_c11 <= Y_15_c10;
               X_16_c11 <= X_16_c10;
               Y_16_c11 <= Y_16_c10;
               X_17_c11 <= X_17_c10;
               Y_17_c11 <= Y_17_c10;
               X_18_c11 <= X_18_c10;
               Y_18_c11 <= Y_18_c10;
               X_19_c11 <= X_19_c10;
               Y_19_c11 <= Y_19_c10;
               X_20_c11 <= X_20_c10;
               Y_20_c11 <= Y_20_c10;
               X_21_c11 <= X_21_c10;
               Y_21_c11 <= Y_21_c10;
               X_22_c11 <= X_22_c10;
               Y_22_c11 <= Y_22_c10;
               X_23_c11 <= X_23_c10;
               Y_23_c11 <= Y_23_c10;
               X_24_c11 <= X_24_c10;
               Y_24_c11 <= Y_24_c10;
               X_25_c11 <= X_25_c10;
               Y_25_c11 <= Y_25_c10;
               X_26_c11 <= X_26_c10;
               Y_26_c11 <= Y_26_c10;
               X_27_c11 <= X_27_c10;
               Y_27_c11 <= Y_27_c10;
            end if;
            if ce_12 = '1' then
               R_0_c12 <= R_0_c11;
               R_1_c12 <= R_1_c11;
               R_2_c12 <= R_2_c11;
               R_3_c12 <= R_3_c11;
               R_4_c12 <= R_4_c11;
               R_5_c12 <= R_5_c11;
               R_6_c12 <= R_6_c11;
               Cin_7_c12 <= Cin_7_c11;
               X_7_c12 <= X_7_c11;
               Y_7_c12 <= Y_7_c11;
               X_8_c12 <= X_8_c11;
               Y_8_c12 <= Y_8_c11;
               X_9_c12 <= X_9_c11;
               Y_9_c12 <= Y_9_c11;
               X_10_c12 <= X_10_c11;
               Y_10_c12 <= Y_10_c11;
               X_11_c12 <= X_11_c11;
               Y_11_c12 <= Y_11_c11;
               X_12_c12 <= X_12_c11;
               Y_12_c12 <= Y_12_c11;
               X_13_c12 <= X_13_c11;
               Y_13_c12 <= Y_13_c11;
               X_14_c12 <= X_14_c11;
               Y_14_c12 <= Y_14_c11;
               X_15_c12 <= X_15_c11;
               Y_15_c12 <= Y_15_c11;
               X_16_c12 <= X_16_c11;
               Y_16_c12 <= Y_16_c11;
               X_17_c12 <= X_17_c11;
               Y_17_c12 <= Y_17_c11;
               X_18_c12 <= X_18_c11;
               Y_18_c12 <= Y_18_c11;
               X_19_c12 <= X_19_c11;
               Y_19_c12 <= Y_19_c11;
               X_20_c12 <= X_20_c11;
               Y_20_c12 <= Y_20_c11;
               X_21_c12 <= X_21_c11;
               Y_21_c12 <= Y_21_c11;
               X_22_c12 <= X_22_c11;
               Y_22_c12 <= Y_22_c11;
               X_23_c12 <= X_23_c11;
               Y_23_c12 <= Y_23_c11;
               X_24_c12 <= X_24_c11;
               Y_24_c12 <= Y_24_c11;
               X_25_c12 <= X_25_c11;
               Y_25_c12 <= Y_25_c11;
               X_26_c12 <= X_26_c11;
               Y_26_c12 <= Y_26_c11;
               X_27_c12 <= X_27_c11;
               Y_27_c12 <= Y_27_c11;
            end if;
            if ce_13 = '1' then
               R_0_c13 <= R_0_c12;
               R_1_c13 <= R_1_c12;
               R_2_c13 <= R_2_c12;
               R_3_c13 <= R_3_c12;
               R_4_c13 <= R_4_c12;
               R_5_c13 <= R_5_c12;
               R_6_c13 <= R_6_c12;
               R_7_c13 <= R_7_c12;
               Cin_8_c13 <= Cin_8_c12;
               X_8_c13 <= X_8_c12;
               Y_8_c13 <= Y_8_c12;
               X_9_c13 <= X_9_c12;
               Y_9_c13 <= Y_9_c12;
               X_10_c13 <= X_10_c12;
               Y_10_c13 <= Y_10_c12;
               X_11_c13 <= X_11_c12;
               Y_11_c13 <= Y_11_c12;
               X_12_c13 <= X_12_c12;
               Y_12_c13 <= Y_12_c12;
               X_13_c13 <= X_13_c12;
               Y_13_c13 <= Y_13_c12;
               X_14_c13 <= X_14_c12;
               Y_14_c13 <= Y_14_c12;
               X_15_c13 <= X_15_c12;
               Y_15_c13 <= Y_15_c12;
               X_16_c13 <= X_16_c12;
               Y_16_c13 <= Y_16_c12;
               X_17_c13 <= X_17_c12;
               Y_17_c13 <= Y_17_c12;
               X_18_c13 <= X_18_c12;
               Y_18_c13 <= Y_18_c12;
               X_19_c13 <= X_19_c12;
               Y_19_c13 <= Y_19_c12;
               X_20_c13 <= X_20_c12;
               Y_20_c13 <= Y_20_c12;
               X_21_c13 <= X_21_c12;
               Y_21_c13 <= Y_21_c12;
               X_22_c13 <= X_22_c12;
               Y_22_c13 <= Y_22_c12;
               X_23_c13 <= X_23_c12;
               Y_23_c13 <= Y_23_c12;
               X_24_c13 <= X_24_c12;
               Y_24_c13 <= Y_24_c12;
               X_25_c13 <= X_25_c12;
               Y_25_c13 <= Y_25_c12;
               X_26_c13 <= X_26_c12;
               Y_26_c13 <= Y_26_c12;
               X_27_c13 <= X_27_c12;
               Y_27_c13 <= Y_27_c12;
            end if;
            if ce_14 = '1' then
               R_0_c14 <= R_0_c13;
               R_1_c14 <= R_1_c13;
               R_2_c14 <= R_2_c13;
               R_3_c14 <= R_3_c13;
               R_4_c14 <= R_4_c13;
               R_5_c14 <= R_5_c13;
               R_6_c14 <= R_6_c13;
               R_7_c14 <= R_7_c13;
               R_8_c14 <= R_8_c13;
               Cin_9_c14 <= Cin_9_c13;
               X_9_c14 <= X_9_c13;
               Y_9_c14 <= Y_9_c13;
               X_10_c14 <= X_10_c13;
               Y_10_c14 <= Y_10_c13;
               X_11_c14 <= X_11_c13;
               Y_11_c14 <= Y_11_c13;
               X_12_c14 <= X_12_c13;
               Y_12_c14 <= Y_12_c13;
               X_13_c14 <= X_13_c13;
               Y_13_c14 <= Y_13_c13;
               X_14_c14 <= X_14_c13;
               Y_14_c14 <= Y_14_c13;
               X_15_c14 <= X_15_c13;
               Y_15_c14 <= Y_15_c13;
               X_16_c14 <= X_16_c13;
               Y_16_c14 <= Y_16_c13;
               X_17_c14 <= X_17_c13;
               Y_17_c14 <= Y_17_c13;
               X_18_c14 <= X_18_c13;
               Y_18_c14 <= Y_18_c13;
               X_19_c14 <= X_19_c13;
               Y_19_c14 <= Y_19_c13;
               X_20_c14 <= X_20_c13;
               Y_20_c14 <= Y_20_c13;
               X_21_c14 <= X_21_c13;
               Y_21_c14 <= Y_21_c13;
               X_22_c14 <= X_22_c13;
               Y_22_c14 <= Y_22_c13;
               X_23_c14 <= X_23_c13;
               Y_23_c14 <= Y_23_c13;
               X_24_c14 <= X_24_c13;
               Y_24_c14 <= Y_24_c13;
               X_25_c14 <= X_25_c13;
               Y_25_c14 <= Y_25_c13;
               X_26_c14 <= X_26_c13;
               Y_26_c14 <= Y_26_c13;
               X_27_c14 <= X_27_c13;
               Y_27_c14 <= Y_27_c13;
            end if;
            if ce_15 = '1' then
               R_0_c15 <= R_0_c14;
               R_1_c15 <= R_1_c14;
               R_2_c15 <= R_2_c14;
               R_3_c15 <= R_3_c14;
               R_4_c15 <= R_4_c14;
               R_5_c15 <= R_5_c14;
               R_6_c15 <= R_6_c14;
               R_7_c15 <= R_7_c14;
               R_8_c15 <= R_8_c14;
               R_9_c15 <= R_9_c14;
               Cin_10_c15 <= Cin_10_c14;
               X_10_c15 <= X_10_c14;
               Y_10_c15 <= Y_10_c14;
               X_11_c15 <= X_11_c14;
               Y_11_c15 <= Y_11_c14;
               X_12_c15 <= X_12_c14;
               Y_12_c15 <= Y_12_c14;
               X_13_c15 <= X_13_c14;
               Y_13_c15 <= Y_13_c14;
               X_14_c15 <= X_14_c14;
               Y_14_c15 <= Y_14_c14;
               X_15_c15 <= X_15_c14;
               Y_15_c15 <= Y_15_c14;
               X_16_c15 <= X_16_c14;
               Y_16_c15 <= Y_16_c14;
               X_17_c15 <= X_17_c14;
               Y_17_c15 <= Y_17_c14;
               X_18_c15 <= X_18_c14;
               Y_18_c15 <= Y_18_c14;
               X_19_c15 <= X_19_c14;
               Y_19_c15 <= Y_19_c14;
               X_20_c15 <= X_20_c14;
               Y_20_c15 <= Y_20_c14;
               X_21_c15 <= X_21_c14;
               Y_21_c15 <= Y_21_c14;
               X_22_c15 <= X_22_c14;
               Y_22_c15 <= Y_22_c14;
               X_23_c15 <= X_23_c14;
               Y_23_c15 <= Y_23_c14;
               X_24_c15 <= X_24_c14;
               Y_24_c15 <= Y_24_c14;
               X_25_c15 <= X_25_c14;
               Y_25_c15 <= Y_25_c14;
               X_26_c15 <= X_26_c14;
               Y_26_c15 <= Y_26_c14;
               X_27_c15 <= X_27_c14;
               Y_27_c15 <= Y_27_c14;
            end if;
            if ce_16 = '1' then
               R_0_c16 <= R_0_c15;
               R_1_c16 <= R_1_c15;
               R_2_c16 <= R_2_c15;
               R_3_c16 <= R_3_c15;
               R_4_c16 <= R_4_c15;
               R_5_c16 <= R_5_c15;
               R_6_c16 <= R_6_c15;
               R_7_c16 <= R_7_c15;
               R_8_c16 <= R_8_c15;
               R_9_c16 <= R_9_c15;
               R_10_c16 <= R_10_c15;
               Cin_11_c16 <= Cin_11_c15;
               X_11_c16 <= X_11_c15;
               Y_11_c16 <= Y_11_c15;
               X_12_c16 <= X_12_c15;
               Y_12_c16 <= Y_12_c15;
               X_13_c16 <= X_13_c15;
               Y_13_c16 <= Y_13_c15;
               X_14_c16 <= X_14_c15;
               Y_14_c16 <= Y_14_c15;
               X_15_c16 <= X_15_c15;
               Y_15_c16 <= Y_15_c15;
               X_16_c16 <= X_16_c15;
               Y_16_c16 <= Y_16_c15;
               X_17_c16 <= X_17_c15;
               Y_17_c16 <= Y_17_c15;
               X_18_c16 <= X_18_c15;
               Y_18_c16 <= Y_18_c15;
               X_19_c16 <= X_19_c15;
               Y_19_c16 <= Y_19_c15;
               X_20_c16 <= X_20_c15;
               Y_20_c16 <= Y_20_c15;
               X_21_c16 <= X_21_c15;
               Y_21_c16 <= Y_21_c15;
               X_22_c16 <= X_22_c15;
               Y_22_c16 <= Y_22_c15;
               X_23_c16 <= X_23_c15;
               Y_23_c16 <= Y_23_c15;
               X_24_c16 <= X_24_c15;
               Y_24_c16 <= Y_24_c15;
               X_25_c16 <= X_25_c15;
               Y_25_c16 <= Y_25_c15;
               X_26_c16 <= X_26_c15;
               Y_26_c16 <= Y_26_c15;
               X_27_c16 <= X_27_c15;
               Y_27_c16 <= Y_27_c15;
            end if;
            if ce_17 = '1' then
               R_0_c17 <= R_0_c16;
               R_1_c17 <= R_1_c16;
               R_2_c17 <= R_2_c16;
               R_3_c17 <= R_3_c16;
               R_4_c17 <= R_4_c16;
               R_5_c17 <= R_5_c16;
               R_6_c17 <= R_6_c16;
               R_7_c17 <= R_7_c16;
               R_8_c17 <= R_8_c16;
               R_9_c17 <= R_9_c16;
               R_10_c17 <= R_10_c16;
               R_11_c17 <= R_11_c16;
               Cin_12_c17 <= Cin_12_c16;
               X_12_c17 <= X_12_c16;
               Y_12_c17 <= Y_12_c16;
               X_13_c17 <= X_13_c16;
               Y_13_c17 <= Y_13_c16;
               X_14_c17 <= X_14_c16;
               Y_14_c17 <= Y_14_c16;
               X_15_c17 <= X_15_c16;
               Y_15_c17 <= Y_15_c16;
               X_16_c17 <= X_16_c16;
               Y_16_c17 <= Y_16_c16;
               X_17_c17 <= X_17_c16;
               Y_17_c17 <= Y_17_c16;
               X_18_c17 <= X_18_c16;
               Y_18_c17 <= Y_18_c16;
               X_19_c17 <= X_19_c16;
               Y_19_c17 <= Y_19_c16;
               X_20_c17 <= X_20_c16;
               Y_20_c17 <= Y_20_c16;
               X_21_c17 <= X_21_c16;
               Y_21_c17 <= Y_21_c16;
               X_22_c17 <= X_22_c16;
               Y_22_c17 <= Y_22_c16;
               X_23_c17 <= X_23_c16;
               Y_23_c17 <= Y_23_c16;
               X_24_c17 <= X_24_c16;
               Y_24_c17 <= Y_24_c16;
               X_25_c17 <= X_25_c16;
               Y_25_c17 <= Y_25_c16;
               X_26_c17 <= X_26_c16;
               Y_26_c17 <= Y_26_c16;
               X_27_c17 <= X_27_c16;
               Y_27_c17 <= Y_27_c16;
            end if;
            if ce_18 = '1' then
               R_0_c18 <= R_0_c17;
               R_1_c18 <= R_1_c17;
               R_2_c18 <= R_2_c17;
               R_3_c18 <= R_3_c17;
               R_4_c18 <= R_4_c17;
               R_5_c18 <= R_5_c17;
               R_6_c18 <= R_6_c17;
               R_7_c18 <= R_7_c17;
               R_8_c18 <= R_8_c17;
               R_9_c18 <= R_9_c17;
               R_10_c18 <= R_10_c17;
               R_11_c18 <= R_11_c17;
               R_12_c18 <= R_12_c17;
               Cin_13_c18 <= Cin_13_c17;
               X_13_c18 <= X_13_c17;
               Y_13_c18 <= Y_13_c17;
               X_14_c18 <= X_14_c17;
               Y_14_c18 <= Y_14_c17;
               X_15_c18 <= X_15_c17;
               Y_15_c18 <= Y_15_c17;
               X_16_c18 <= X_16_c17;
               Y_16_c18 <= Y_16_c17;
               X_17_c18 <= X_17_c17;
               Y_17_c18 <= Y_17_c17;
               X_18_c18 <= X_18_c17;
               Y_18_c18 <= Y_18_c17;
               X_19_c18 <= X_19_c17;
               Y_19_c18 <= Y_19_c17;
               X_20_c18 <= X_20_c17;
               Y_20_c18 <= Y_20_c17;
               X_21_c18 <= X_21_c17;
               Y_21_c18 <= Y_21_c17;
               X_22_c18 <= X_22_c17;
               Y_22_c18 <= Y_22_c17;
               X_23_c18 <= X_23_c17;
               Y_23_c18 <= Y_23_c17;
               X_24_c18 <= X_24_c17;
               Y_24_c18 <= Y_24_c17;
               X_25_c18 <= X_25_c17;
               Y_25_c18 <= Y_25_c17;
               X_26_c18 <= X_26_c17;
               Y_26_c18 <= Y_26_c17;
               X_27_c18 <= X_27_c17;
               Y_27_c18 <= Y_27_c17;
            end if;
            if ce_19 = '1' then
               R_0_c19 <= R_0_c18;
               R_1_c19 <= R_1_c18;
               R_2_c19 <= R_2_c18;
               R_3_c19 <= R_3_c18;
               R_4_c19 <= R_4_c18;
               R_5_c19 <= R_5_c18;
               R_6_c19 <= R_6_c18;
               R_7_c19 <= R_7_c18;
               R_8_c19 <= R_8_c18;
               R_9_c19 <= R_9_c18;
               R_10_c19 <= R_10_c18;
               R_11_c19 <= R_11_c18;
               R_12_c19 <= R_12_c18;
               R_13_c19 <= R_13_c18;
               Cin_14_c19 <= Cin_14_c18;
               X_14_c19 <= X_14_c18;
               Y_14_c19 <= Y_14_c18;
               X_15_c19 <= X_15_c18;
               Y_15_c19 <= Y_15_c18;
               X_16_c19 <= X_16_c18;
               Y_16_c19 <= Y_16_c18;
               X_17_c19 <= X_17_c18;
               Y_17_c19 <= Y_17_c18;
               X_18_c19 <= X_18_c18;
               Y_18_c19 <= Y_18_c18;
               X_19_c19 <= X_19_c18;
               Y_19_c19 <= Y_19_c18;
               X_20_c19 <= X_20_c18;
               Y_20_c19 <= Y_20_c18;
               X_21_c19 <= X_21_c18;
               Y_21_c19 <= Y_21_c18;
               X_22_c19 <= X_22_c18;
               Y_22_c19 <= Y_22_c18;
               X_23_c19 <= X_23_c18;
               Y_23_c19 <= Y_23_c18;
               X_24_c19 <= X_24_c18;
               Y_24_c19 <= Y_24_c18;
               X_25_c19 <= X_25_c18;
               Y_25_c19 <= Y_25_c18;
               X_26_c19 <= X_26_c18;
               Y_26_c19 <= Y_26_c18;
               X_27_c19 <= X_27_c18;
               Y_27_c19 <= Y_27_c18;
            end if;
            if ce_20 = '1' then
               R_0_c20 <= R_0_c19;
               R_1_c20 <= R_1_c19;
               R_2_c20 <= R_2_c19;
               R_3_c20 <= R_3_c19;
               R_4_c20 <= R_4_c19;
               R_5_c20 <= R_5_c19;
               R_6_c20 <= R_6_c19;
               R_7_c20 <= R_7_c19;
               R_8_c20 <= R_8_c19;
               R_9_c20 <= R_9_c19;
               R_10_c20 <= R_10_c19;
               R_11_c20 <= R_11_c19;
               R_12_c20 <= R_12_c19;
               R_13_c20 <= R_13_c19;
               Cin_14_c20 <= Cin_14_c19;
               X_14_c20 <= X_14_c19;
               Y_14_c20 <= Y_14_c19;
               X_15_c20 <= X_15_c19;
               Y_15_c20 <= Y_15_c19;
               X_16_c20 <= X_16_c19;
               Y_16_c20 <= Y_16_c19;
               X_17_c20 <= X_17_c19;
               Y_17_c20 <= Y_17_c19;
               X_18_c20 <= X_18_c19;
               Y_18_c20 <= Y_18_c19;
               X_19_c20 <= X_19_c19;
               Y_19_c20 <= Y_19_c19;
               X_20_c20 <= X_20_c19;
               Y_20_c20 <= Y_20_c19;
               X_21_c20 <= X_21_c19;
               Y_21_c20 <= Y_21_c19;
               X_22_c20 <= X_22_c19;
               Y_22_c20 <= Y_22_c19;
               X_23_c20 <= X_23_c19;
               Y_23_c20 <= Y_23_c19;
               X_24_c20 <= X_24_c19;
               Y_24_c20 <= Y_24_c19;
               X_25_c20 <= X_25_c19;
               Y_25_c20 <= Y_25_c19;
               X_26_c20 <= X_26_c19;
               Y_26_c20 <= Y_26_c19;
               X_27_c20 <= X_27_c19;
               Y_27_c20 <= Y_27_c19;
            end if;
            if ce_21 = '1' then
               R_0_c21 <= R_0_c20;
               R_1_c21 <= R_1_c20;
               R_2_c21 <= R_2_c20;
               R_3_c21 <= R_3_c20;
               R_4_c21 <= R_4_c20;
               R_5_c21 <= R_5_c20;
               R_6_c21 <= R_6_c20;
               R_7_c21 <= R_7_c20;
               R_8_c21 <= R_8_c20;
               R_9_c21 <= R_9_c20;
               R_10_c21 <= R_10_c20;
               R_11_c21 <= R_11_c20;
               R_12_c21 <= R_12_c20;
               R_13_c21 <= R_13_c20;
               R_14_c21 <= R_14_c20;
               Cin_15_c21 <= Cin_15_c20;
               X_15_c21 <= X_15_c20;
               Y_15_c21 <= Y_15_c20;
               X_16_c21 <= X_16_c20;
               Y_16_c21 <= Y_16_c20;
               X_17_c21 <= X_17_c20;
               Y_17_c21 <= Y_17_c20;
               X_18_c21 <= X_18_c20;
               Y_18_c21 <= Y_18_c20;
               X_19_c21 <= X_19_c20;
               Y_19_c21 <= Y_19_c20;
               X_20_c21 <= X_20_c20;
               Y_20_c21 <= Y_20_c20;
               X_21_c21 <= X_21_c20;
               Y_21_c21 <= Y_21_c20;
               X_22_c21 <= X_22_c20;
               Y_22_c21 <= Y_22_c20;
               X_23_c21 <= X_23_c20;
               Y_23_c21 <= Y_23_c20;
               X_24_c21 <= X_24_c20;
               Y_24_c21 <= Y_24_c20;
               X_25_c21 <= X_25_c20;
               Y_25_c21 <= Y_25_c20;
               X_26_c21 <= X_26_c20;
               Y_26_c21 <= Y_26_c20;
               X_27_c21 <= X_27_c20;
               Y_27_c21 <= Y_27_c20;
            end if;
            if ce_22 = '1' then
               R_0_c22 <= R_0_c21;
               R_1_c22 <= R_1_c21;
               R_2_c22 <= R_2_c21;
               R_3_c22 <= R_3_c21;
               R_4_c22 <= R_4_c21;
               R_5_c22 <= R_5_c21;
               R_6_c22 <= R_6_c21;
               R_7_c22 <= R_7_c21;
               R_8_c22 <= R_8_c21;
               R_9_c22 <= R_9_c21;
               R_10_c22 <= R_10_c21;
               R_11_c22 <= R_11_c21;
               R_12_c22 <= R_12_c21;
               R_13_c22 <= R_13_c21;
               R_14_c22 <= R_14_c21;
               R_15_c22 <= R_15_c21;
               Cin_16_c22 <= Cin_16_c21;
               X_16_c22 <= X_16_c21;
               Y_16_c22 <= Y_16_c21;
               X_17_c22 <= X_17_c21;
               Y_17_c22 <= Y_17_c21;
               X_18_c22 <= X_18_c21;
               Y_18_c22 <= Y_18_c21;
               X_19_c22 <= X_19_c21;
               Y_19_c22 <= Y_19_c21;
               X_20_c22 <= X_20_c21;
               Y_20_c22 <= Y_20_c21;
               X_21_c22 <= X_21_c21;
               Y_21_c22 <= Y_21_c21;
               X_22_c22 <= X_22_c21;
               Y_22_c22 <= Y_22_c21;
               X_23_c22 <= X_23_c21;
               Y_23_c22 <= Y_23_c21;
               X_24_c22 <= X_24_c21;
               Y_24_c22 <= Y_24_c21;
               X_25_c22 <= X_25_c21;
               Y_25_c22 <= Y_25_c21;
               X_26_c22 <= X_26_c21;
               Y_26_c22 <= Y_26_c21;
               X_27_c22 <= X_27_c21;
               Y_27_c22 <= Y_27_c21;
            end if;
            if ce_23 = '1' then
               R_0_c23 <= R_0_c22;
               R_1_c23 <= R_1_c22;
               R_2_c23 <= R_2_c22;
               R_3_c23 <= R_3_c22;
               R_4_c23 <= R_4_c22;
               R_5_c23 <= R_5_c22;
               R_6_c23 <= R_6_c22;
               R_7_c23 <= R_7_c22;
               R_8_c23 <= R_8_c22;
               R_9_c23 <= R_9_c22;
               R_10_c23 <= R_10_c22;
               R_11_c23 <= R_11_c22;
               R_12_c23 <= R_12_c22;
               R_13_c23 <= R_13_c22;
               R_14_c23 <= R_14_c22;
               R_15_c23 <= R_15_c22;
               R_16_c23 <= R_16_c22;
               Cin_17_c23 <= Cin_17_c22;
               X_17_c23 <= X_17_c22;
               Y_17_c23 <= Y_17_c22;
               X_18_c23 <= X_18_c22;
               Y_18_c23 <= Y_18_c22;
               X_19_c23 <= X_19_c22;
               Y_19_c23 <= Y_19_c22;
               X_20_c23 <= X_20_c22;
               Y_20_c23 <= Y_20_c22;
               X_21_c23 <= X_21_c22;
               Y_21_c23 <= Y_21_c22;
               X_22_c23 <= X_22_c22;
               Y_22_c23 <= Y_22_c22;
               X_23_c23 <= X_23_c22;
               Y_23_c23 <= Y_23_c22;
               X_24_c23 <= X_24_c22;
               Y_24_c23 <= Y_24_c22;
               X_25_c23 <= X_25_c22;
               Y_25_c23 <= Y_25_c22;
               X_26_c23 <= X_26_c22;
               Y_26_c23 <= Y_26_c22;
               X_27_c23 <= X_27_c22;
               Y_27_c23 <= Y_27_c22;
            end if;
            if ce_24 = '1' then
               R_0_c24 <= R_0_c23;
               R_1_c24 <= R_1_c23;
               R_2_c24 <= R_2_c23;
               R_3_c24 <= R_3_c23;
               R_4_c24 <= R_4_c23;
               R_5_c24 <= R_5_c23;
               R_6_c24 <= R_6_c23;
               R_7_c24 <= R_7_c23;
               R_8_c24 <= R_8_c23;
               R_9_c24 <= R_9_c23;
               R_10_c24 <= R_10_c23;
               R_11_c24 <= R_11_c23;
               R_12_c24 <= R_12_c23;
               R_13_c24 <= R_13_c23;
               R_14_c24 <= R_14_c23;
               R_15_c24 <= R_15_c23;
               R_16_c24 <= R_16_c23;
               R_17_c24 <= R_17_c23;
               Cin_18_c24 <= Cin_18_c23;
               X_18_c24 <= X_18_c23;
               Y_18_c24 <= Y_18_c23;
               X_19_c24 <= X_19_c23;
               Y_19_c24 <= Y_19_c23;
               X_20_c24 <= X_20_c23;
               Y_20_c24 <= Y_20_c23;
               X_21_c24 <= X_21_c23;
               Y_21_c24 <= Y_21_c23;
               X_22_c24 <= X_22_c23;
               Y_22_c24 <= Y_22_c23;
               X_23_c24 <= X_23_c23;
               Y_23_c24 <= Y_23_c23;
               X_24_c24 <= X_24_c23;
               Y_24_c24 <= Y_24_c23;
               X_25_c24 <= X_25_c23;
               Y_25_c24 <= Y_25_c23;
               X_26_c24 <= X_26_c23;
               Y_26_c24 <= Y_26_c23;
               X_27_c24 <= X_27_c23;
               Y_27_c24 <= Y_27_c23;
            end if;
            if ce_25 = '1' then
               R_0_c25 <= R_0_c24;
               R_1_c25 <= R_1_c24;
               R_2_c25 <= R_2_c24;
               R_3_c25 <= R_3_c24;
               R_4_c25 <= R_4_c24;
               R_5_c25 <= R_5_c24;
               R_6_c25 <= R_6_c24;
               R_7_c25 <= R_7_c24;
               R_8_c25 <= R_8_c24;
               R_9_c25 <= R_9_c24;
               R_10_c25 <= R_10_c24;
               R_11_c25 <= R_11_c24;
               R_12_c25 <= R_12_c24;
               R_13_c25 <= R_13_c24;
               R_14_c25 <= R_14_c24;
               R_15_c25 <= R_15_c24;
               R_16_c25 <= R_16_c24;
               R_17_c25 <= R_17_c24;
               R_18_c25 <= R_18_c24;
               Cin_19_c25 <= Cin_19_c24;
               X_19_c25 <= X_19_c24;
               Y_19_c25 <= Y_19_c24;
               X_20_c25 <= X_20_c24;
               Y_20_c25 <= Y_20_c24;
               X_21_c25 <= X_21_c24;
               Y_21_c25 <= Y_21_c24;
               X_22_c25 <= X_22_c24;
               Y_22_c25 <= Y_22_c24;
               X_23_c25 <= X_23_c24;
               Y_23_c25 <= Y_23_c24;
               X_24_c25 <= X_24_c24;
               Y_24_c25 <= Y_24_c24;
               X_25_c25 <= X_25_c24;
               Y_25_c25 <= Y_25_c24;
               X_26_c25 <= X_26_c24;
               Y_26_c25 <= Y_26_c24;
               X_27_c25 <= X_27_c24;
               Y_27_c25 <= Y_27_c24;
            end if;
            if ce_26 = '1' then
               R_0_c26 <= R_0_c25;
               R_1_c26 <= R_1_c25;
               R_2_c26 <= R_2_c25;
               R_3_c26 <= R_3_c25;
               R_4_c26 <= R_4_c25;
               R_5_c26 <= R_5_c25;
               R_6_c26 <= R_6_c25;
               R_7_c26 <= R_7_c25;
               R_8_c26 <= R_8_c25;
               R_9_c26 <= R_9_c25;
               R_10_c26 <= R_10_c25;
               R_11_c26 <= R_11_c25;
               R_12_c26 <= R_12_c25;
               R_13_c26 <= R_13_c25;
               R_14_c26 <= R_14_c25;
               R_15_c26 <= R_15_c25;
               R_16_c26 <= R_16_c25;
               R_17_c26 <= R_17_c25;
               R_18_c26 <= R_18_c25;
               R_19_c26 <= R_19_c25;
               Cin_20_c26 <= Cin_20_c25;
               X_20_c26 <= X_20_c25;
               Y_20_c26 <= Y_20_c25;
               X_21_c26 <= X_21_c25;
               Y_21_c26 <= Y_21_c25;
               X_22_c26 <= X_22_c25;
               Y_22_c26 <= Y_22_c25;
               X_23_c26 <= X_23_c25;
               Y_23_c26 <= Y_23_c25;
               X_24_c26 <= X_24_c25;
               Y_24_c26 <= Y_24_c25;
               X_25_c26 <= X_25_c25;
               Y_25_c26 <= Y_25_c25;
               X_26_c26 <= X_26_c25;
               Y_26_c26 <= Y_26_c25;
               X_27_c26 <= X_27_c25;
               Y_27_c26 <= Y_27_c25;
            end if;
            if ce_27 = '1' then
               R_0_c27 <= R_0_c26;
               R_1_c27 <= R_1_c26;
               R_2_c27 <= R_2_c26;
               R_3_c27 <= R_3_c26;
               R_4_c27 <= R_4_c26;
               R_5_c27 <= R_5_c26;
               R_6_c27 <= R_6_c26;
               R_7_c27 <= R_7_c26;
               R_8_c27 <= R_8_c26;
               R_9_c27 <= R_9_c26;
               R_10_c27 <= R_10_c26;
               R_11_c27 <= R_11_c26;
               R_12_c27 <= R_12_c26;
               R_13_c27 <= R_13_c26;
               R_14_c27 <= R_14_c26;
               R_15_c27 <= R_15_c26;
               R_16_c27 <= R_16_c26;
               R_17_c27 <= R_17_c26;
               R_18_c27 <= R_18_c26;
               R_19_c27 <= R_19_c26;
               R_20_c27 <= R_20_c26;
               Cin_21_c27 <= Cin_21_c26;
               X_21_c27 <= X_21_c26;
               Y_21_c27 <= Y_21_c26;
               X_22_c27 <= X_22_c26;
               Y_22_c27 <= Y_22_c26;
               X_23_c27 <= X_23_c26;
               Y_23_c27 <= Y_23_c26;
               X_24_c27 <= X_24_c26;
               Y_24_c27 <= Y_24_c26;
               X_25_c27 <= X_25_c26;
               Y_25_c27 <= Y_25_c26;
               X_26_c27 <= X_26_c26;
               Y_26_c27 <= Y_26_c26;
               X_27_c27 <= X_27_c26;
               Y_27_c27 <= Y_27_c26;
            end if;
            if ce_28 = '1' then
               R_0_c28 <= R_0_c27;
               R_1_c28 <= R_1_c27;
               R_2_c28 <= R_2_c27;
               R_3_c28 <= R_3_c27;
               R_4_c28 <= R_4_c27;
               R_5_c28 <= R_5_c27;
               R_6_c28 <= R_6_c27;
               R_7_c28 <= R_7_c27;
               R_8_c28 <= R_8_c27;
               R_9_c28 <= R_9_c27;
               R_10_c28 <= R_10_c27;
               R_11_c28 <= R_11_c27;
               R_12_c28 <= R_12_c27;
               R_13_c28 <= R_13_c27;
               R_14_c28 <= R_14_c27;
               R_15_c28 <= R_15_c27;
               R_16_c28 <= R_16_c27;
               R_17_c28 <= R_17_c27;
               R_18_c28 <= R_18_c27;
               R_19_c28 <= R_19_c27;
               R_20_c28 <= R_20_c27;
               R_21_c28 <= R_21_c27;
               Cin_22_c28 <= Cin_22_c27;
               X_22_c28 <= X_22_c27;
               Y_22_c28 <= Y_22_c27;
               X_23_c28 <= X_23_c27;
               Y_23_c28 <= Y_23_c27;
               X_24_c28 <= X_24_c27;
               Y_24_c28 <= Y_24_c27;
               X_25_c28 <= X_25_c27;
               Y_25_c28 <= Y_25_c27;
               X_26_c28 <= X_26_c27;
               Y_26_c28 <= Y_26_c27;
               X_27_c28 <= X_27_c27;
               Y_27_c28 <= Y_27_c27;
            end if;
            if ce_29 = '1' then
               R_0_c29 <= R_0_c28;
               R_1_c29 <= R_1_c28;
               R_2_c29 <= R_2_c28;
               R_3_c29 <= R_3_c28;
               R_4_c29 <= R_4_c28;
               R_5_c29 <= R_5_c28;
               R_6_c29 <= R_6_c28;
               R_7_c29 <= R_7_c28;
               R_8_c29 <= R_8_c28;
               R_9_c29 <= R_9_c28;
               R_10_c29 <= R_10_c28;
               R_11_c29 <= R_11_c28;
               R_12_c29 <= R_12_c28;
               R_13_c29 <= R_13_c28;
               R_14_c29 <= R_14_c28;
               R_15_c29 <= R_15_c28;
               R_16_c29 <= R_16_c28;
               R_17_c29 <= R_17_c28;
               R_18_c29 <= R_18_c28;
               R_19_c29 <= R_19_c28;
               R_20_c29 <= R_20_c28;
               R_21_c29 <= R_21_c28;
               R_22_c29 <= R_22_c28;
               Cin_23_c29 <= Cin_23_c28;
               X_23_c29 <= X_23_c28;
               Y_23_c29 <= Y_23_c28;
               X_24_c29 <= X_24_c28;
               Y_24_c29 <= Y_24_c28;
               X_25_c29 <= X_25_c28;
               Y_25_c29 <= Y_25_c28;
               X_26_c29 <= X_26_c28;
               Y_26_c29 <= Y_26_c28;
               X_27_c29 <= X_27_c28;
               Y_27_c29 <= Y_27_c28;
            end if;
            if ce_30 = '1' then
               R_0_c30 <= R_0_c29;
               R_1_c30 <= R_1_c29;
               R_2_c30 <= R_2_c29;
               R_3_c30 <= R_3_c29;
               R_4_c30 <= R_4_c29;
               R_5_c30 <= R_5_c29;
               R_6_c30 <= R_6_c29;
               R_7_c30 <= R_7_c29;
               R_8_c30 <= R_8_c29;
               R_9_c30 <= R_9_c29;
               R_10_c30 <= R_10_c29;
               R_11_c30 <= R_11_c29;
               R_12_c30 <= R_12_c29;
               R_13_c30 <= R_13_c29;
               R_14_c30 <= R_14_c29;
               R_15_c30 <= R_15_c29;
               R_16_c30 <= R_16_c29;
               R_17_c30 <= R_17_c29;
               R_18_c30 <= R_18_c29;
               R_19_c30 <= R_19_c29;
               R_20_c30 <= R_20_c29;
               R_21_c30 <= R_21_c29;
               R_22_c30 <= R_22_c29;
               R_23_c30 <= R_23_c29;
               Cin_24_c30 <= Cin_24_c29;
               X_24_c30 <= X_24_c29;
               Y_24_c30 <= Y_24_c29;
               X_25_c30 <= X_25_c29;
               Y_25_c30 <= Y_25_c29;
               X_26_c30 <= X_26_c29;
               Y_26_c30 <= Y_26_c29;
               X_27_c30 <= X_27_c29;
               Y_27_c30 <= Y_27_c29;
            end if;
            if ce_31 = '1' then
               R_0_c31 <= R_0_c30;
               R_1_c31 <= R_1_c30;
               R_2_c31 <= R_2_c30;
               R_3_c31 <= R_3_c30;
               R_4_c31 <= R_4_c30;
               R_5_c31 <= R_5_c30;
               R_6_c31 <= R_6_c30;
               R_7_c31 <= R_7_c30;
               R_8_c31 <= R_8_c30;
               R_9_c31 <= R_9_c30;
               R_10_c31 <= R_10_c30;
               R_11_c31 <= R_11_c30;
               R_12_c31 <= R_12_c30;
               R_13_c31 <= R_13_c30;
               R_14_c31 <= R_14_c30;
               R_15_c31 <= R_15_c30;
               R_16_c31 <= R_16_c30;
               R_17_c31 <= R_17_c30;
               R_18_c31 <= R_18_c30;
               R_19_c31 <= R_19_c30;
               R_20_c31 <= R_20_c30;
               R_21_c31 <= R_21_c30;
               R_22_c31 <= R_22_c30;
               R_23_c31 <= R_23_c30;
               R_24_c31 <= R_24_c30;
               Cin_25_c31 <= Cin_25_c30;
               X_25_c31 <= X_25_c30;
               Y_25_c31 <= Y_25_c30;
               X_26_c31 <= X_26_c30;
               Y_26_c31 <= Y_26_c30;
               X_27_c31 <= X_27_c30;
               Y_27_c31 <= Y_27_c30;
            end if;
            if ce_32 = '1' then
               R_0_c32 <= R_0_c31;
               R_1_c32 <= R_1_c31;
               R_2_c32 <= R_2_c31;
               R_3_c32 <= R_3_c31;
               R_4_c32 <= R_4_c31;
               R_5_c32 <= R_5_c31;
               R_6_c32 <= R_6_c31;
               R_7_c32 <= R_7_c31;
               R_8_c32 <= R_8_c31;
               R_9_c32 <= R_9_c31;
               R_10_c32 <= R_10_c31;
               R_11_c32 <= R_11_c31;
               R_12_c32 <= R_12_c31;
               R_13_c32 <= R_13_c31;
               R_14_c32 <= R_14_c31;
               R_15_c32 <= R_15_c31;
               R_16_c32 <= R_16_c31;
               R_17_c32 <= R_17_c31;
               R_18_c32 <= R_18_c31;
               R_19_c32 <= R_19_c31;
               R_20_c32 <= R_20_c31;
               R_21_c32 <= R_21_c31;
               R_22_c32 <= R_22_c31;
               R_23_c32 <= R_23_c31;
               R_24_c32 <= R_24_c31;
               R_25_c32 <= R_25_c31;
               Cin_26_c32 <= Cin_26_c31;
               X_26_c32 <= X_26_c31;
               Y_26_c32 <= Y_26_c31;
               X_27_c32 <= X_27_c31;
               Y_27_c32 <= Y_27_c31;
            end if;
            if ce_33 = '1' then
               R_0_c33 <= R_0_c32;
               R_1_c33 <= R_1_c32;
               R_2_c33 <= R_2_c32;
               R_3_c33 <= R_3_c32;
               R_4_c33 <= R_4_c32;
               R_5_c33 <= R_5_c32;
               R_6_c33 <= R_6_c32;
               R_7_c33 <= R_7_c32;
               R_8_c33 <= R_8_c32;
               R_9_c33 <= R_9_c32;
               R_10_c33 <= R_10_c32;
               R_11_c33 <= R_11_c32;
               R_12_c33 <= R_12_c32;
               R_13_c33 <= R_13_c32;
               R_14_c33 <= R_14_c32;
               R_15_c33 <= R_15_c32;
               R_16_c33 <= R_16_c32;
               R_17_c33 <= R_17_c32;
               R_18_c33 <= R_18_c32;
               R_19_c33 <= R_19_c32;
               R_20_c33 <= R_20_c32;
               R_21_c33 <= R_21_c32;
               R_22_c33 <= R_22_c32;
               R_23_c33 <= R_23_c32;
               R_24_c33 <= R_24_c32;
               R_25_c33 <= R_25_c32;
               R_26_c33 <= R_26_c32;
               Cin_27_c33 <= Cin_27_c32;
               X_27_c33 <= X_27_c32;
               Y_27_c33 <= Y_27_c32;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c4 <= '0' & X(2 downto 0);
   Y_0_c4 <= '0' & Y(2 downto 0);
   S_0_c5 <= X_0_c5 + Y_0_c5 + Cin_0_c5;
   R_0_c5 <= S_0_c5(2 downto 0);
   Cin_1_c5 <= S_0_c5(3);
   X_1_c4 <= '0' & X(5 downto 3);
   Y_1_c4 <= '0' & Y(5 downto 3);
   S_1_c6 <= X_1_c6 + Y_1_c6 + Cin_1_c6;
   R_1_c6 <= S_1_c6(2 downto 0);
   Cin_2_c6 <= S_1_c6(3);
   X_2_c4 <= '0' & X(8 downto 6);
   Y_2_c4 <= '0' & Y(8 downto 6);
   S_2_c7 <= X_2_c7 + Y_2_c7 + Cin_2_c7;
   R_2_c7 <= S_2_c7(2 downto 0);
   Cin_3_c7 <= S_2_c7(3);
   X_3_c4 <= '0' & X(11 downto 9);
   Y_3_c4 <= '0' & Y(11 downto 9);
   S_3_c8 <= X_3_c8 + Y_3_c8 + Cin_3_c8;
   R_3_c8 <= S_3_c8(2 downto 0);
   Cin_4_c8 <= S_3_c8(3);
   X_4_c4 <= '0' & X(14 downto 12);
   Y_4_c4 <= '0' & Y(14 downto 12);
   S_4_c9 <= X_4_c9 + Y_4_c9 + Cin_4_c9;
   R_4_c9 <= S_4_c9(2 downto 0);
   Cin_5_c9 <= S_4_c9(3);
   X_5_c4 <= '0' & X(17 downto 15);
   Y_5_c4 <= '0' & Y(17 downto 15);
   S_5_c10 <= X_5_c10 + Y_5_c10 + Cin_5_c10;
   R_5_c10 <= S_5_c10(2 downto 0);
   Cin_6_c10 <= S_5_c10(3);
   X_6_c4 <= '0' & X(20 downto 18);
   Y_6_c4 <= '0' & Y(20 downto 18);
   S_6_c11 <= X_6_c11 + Y_6_c11 + Cin_6_c11;
   R_6_c11 <= S_6_c11(2 downto 0);
   Cin_7_c11 <= S_6_c11(3);
   X_7_c4 <= '0' & X(23 downto 21);
   Y_7_c4 <= '0' & Y(23 downto 21);
   S_7_c12 <= X_7_c12 + Y_7_c12 + Cin_7_c12;
   R_7_c12 <= S_7_c12(2 downto 0);
   Cin_8_c12 <= S_7_c12(3);
   X_8_c4 <= '0' & X(26 downto 24);
   Y_8_c4 <= '0' & Y(26 downto 24);
   S_8_c13 <= X_8_c13 + Y_8_c13 + Cin_8_c13;
   R_8_c13 <= S_8_c13(2 downto 0);
   Cin_9_c13 <= S_8_c13(3);
   X_9_c4 <= '0' & X(29 downto 27);
   Y_9_c4 <= '0' & Y(29 downto 27);
   S_9_c14 <= X_9_c14 + Y_9_c14 + Cin_9_c14;
   R_9_c14 <= S_9_c14(2 downto 0);
   Cin_10_c14 <= S_9_c14(3);
   X_10_c4 <= '0' & X(32 downto 30);
   Y_10_c4 <= '0' & Y(32 downto 30);
   S_10_c15 <= X_10_c15 + Y_10_c15 + Cin_10_c15;
   R_10_c15 <= S_10_c15(2 downto 0);
   Cin_11_c15 <= S_10_c15(3);
   X_11_c4 <= '0' & X(35 downto 33);
   Y_11_c4 <= '0' & Y(35 downto 33);
   S_11_c16 <= X_11_c16 + Y_11_c16 + Cin_11_c16;
   R_11_c16 <= S_11_c16(2 downto 0);
   Cin_12_c16 <= S_11_c16(3);
   X_12_c4 <= '0' & X(38 downto 36);
   Y_12_c4 <= '0' & Y(38 downto 36);
   S_12_c17 <= X_12_c17 + Y_12_c17 + Cin_12_c17;
   R_12_c17 <= S_12_c17(2 downto 0);
   Cin_13_c17 <= S_12_c17(3);
   X_13_c4 <= '0' & X(41 downto 39);
   Y_13_c4 <= '0' & Y(41 downto 39);
   S_13_c18 <= X_13_c18 + Y_13_c18 + Cin_13_c18;
   R_13_c18 <= S_13_c18(2 downto 0);
   Cin_14_c18 <= S_13_c18(3);
   X_14_c4 <= '0' & X(44 downto 42);
   Y_14_c4 <= '0' & Y(44 downto 42);
   S_14_c20 <= X_14_c20 + Y_14_c20 + Cin_14_c20;
   R_14_c20 <= S_14_c20(2 downto 0);
   Cin_15_c20 <= S_14_c20(3);
   X_15_c4 <= '0' & X(47 downto 45);
   Y_15_c4 <= '0' & Y(47 downto 45);
   S_15_c21 <= X_15_c21 + Y_15_c21 + Cin_15_c21;
   R_15_c21 <= S_15_c21(2 downto 0);
   Cin_16_c21 <= S_15_c21(3);
   X_16_c4 <= '0' & X(50 downto 48);
   Y_16_c4 <= '0' & Y(50 downto 48);
   S_16_c22 <= X_16_c22 + Y_16_c22 + Cin_16_c22;
   R_16_c22 <= S_16_c22(2 downto 0);
   Cin_17_c22 <= S_16_c22(3);
   X_17_c4 <= '0' & X(53 downto 51);
   Y_17_c4 <= '0' & Y(53 downto 51);
   S_17_c23 <= X_17_c23 + Y_17_c23 + Cin_17_c23;
   R_17_c23 <= S_17_c23(2 downto 0);
   Cin_18_c23 <= S_17_c23(3);
   X_18_c4 <= '0' & X(56 downto 54);
   Y_18_c4 <= '0' & Y(56 downto 54);
   S_18_c24 <= X_18_c24 + Y_18_c24 + Cin_18_c24;
   R_18_c24 <= S_18_c24(2 downto 0);
   Cin_19_c24 <= S_18_c24(3);
   X_19_c4 <= '0' & X(59 downto 57);
   Y_19_c4 <= '0' & Y(59 downto 57);
   S_19_c25 <= X_19_c25 + Y_19_c25 + Cin_19_c25;
   R_19_c25 <= S_19_c25(2 downto 0);
   Cin_20_c25 <= S_19_c25(3);
   X_20_c4 <= '0' & X(62 downto 60);
   Y_20_c4 <= '0' & Y(62 downto 60);
   S_20_c26 <= X_20_c26 + Y_20_c26 + Cin_20_c26;
   R_20_c26 <= S_20_c26(2 downto 0);
   Cin_21_c26 <= S_20_c26(3);
   X_21_c4 <= '0' & X(65 downto 63);
   Y_21_c4 <= '0' & Y(65 downto 63);
   S_21_c27 <= X_21_c27 + Y_21_c27 + Cin_21_c27;
   R_21_c27 <= S_21_c27(2 downto 0);
   Cin_22_c27 <= S_21_c27(3);
   X_22_c4 <= '0' & X(68 downto 66);
   Y_22_c4 <= '0' & Y(68 downto 66);
   S_22_c28 <= X_22_c28 + Y_22_c28 + Cin_22_c28;
   R_22_c28 <= S_22_c28(2 downto 0);
   Cin_23_c28 <= S_22_c28(3);
   X_23_c4 <= '0' & X(71 downto 69);
   Y_23_c4 <= '0' & Y(71 downto 69);
   S_23_c29 <= X_23_c29 + Y_23_c29 + Cin_23_c29;
   R_23_c29 <= S_23_c29(2 downto 0);
   Cin_24_c29 <= S_23_c29(3);
   X_24_c4 <= '0' & X(74 downto 72);
   Y_24_c4 <= '0' & Y(74 downto 72);
   S_24_c30 <= X_24_c30 + Y_24_c30 + Cin_24_c30;
   R_24_c30 <= S_24_c30(2 downto 0);
   Cin_25_c30 <= S_24_c30(3);
   X_25_c4 <= '0' & X(77 downto 75);
   Y_25_c4 <= '0' & Y(77 downto 75);
   S_25_c31 <= X_25_c31 + Y_25_c31 + Cin_25_c31;
   R_25_c31 <= S_25_c31(2 downto 0);
   Cin_26_c31 <= S_25_c31(3);
   X_26_c4 <= '0' & X(80 downto 78);
   Y_26_c4 <= '0' & Y(80 downto 78);
   S_26_c32 <= X_26_c32 + Y_26_c32 + Cin_26_c32;
   R_26_c32 <= S_26_c32(2 downto 0);
   Cin_27_c32 <= S_26_c32(3);
   X_27_c4 <= '0' & X(83 downto 81);
   Y_27_c4 <= '0' & Y(83 downto 81);
   S_27_c33 <= X_27_c33 + Y_27_c33 + Cin_27_c33;
   R_27_c33 <= S_27_c33(2 downto 0);
   R <= R_27_c33 & R_26_c33 & R_25_c33 & R_24_c33 & R_23_c33 & R_22_c33 & R_21_c33 & R_20_c33 & R_19_c33 & R_18_c33 & R_17_c33 & R_16_c33 & R_15_c33 & R_14_c33 & R_13_c33 & R_12_c33 & R_11_c33 & R_10_c33 & R_9_c33 & R_8_c33 & R_7_c33 & R_6_c33 & R_5_c33 & R_4_c33 & R_3_c33 & R_2_c33 & R_1_c33 & R_0_c33 ;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_53x53_106_Freq800_uid5
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_53x53_106_Freq800_uid5 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of IntMultiplier_53x53_106_Freq800_uid5 is
   component DSPBlock_17x24_Freq800_uid9 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid11 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid13 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid40 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid55 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid57 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid59 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid76 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid81 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid86 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid91 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid96 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid101 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid103 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid105 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid111 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid116 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid136 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid141 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid146 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid151 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid156 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid161 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid166 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid171 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid173 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid175 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid177 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid179 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid181 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid191 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid196 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid201 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid206 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid211 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid216 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid221 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid226 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid231 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid236 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid241 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid243 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid245 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid247 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid249 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid251 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid256 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid261 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid266 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid271 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid276 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid281 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid286 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid291 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid296 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid301 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid306 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid311 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid316 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq800_uid322 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq800_uid326 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq800_uid334 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq800_uid400 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq800_uid432 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntAdder_84_Freq800_uid972 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
             X : in  std_logic_vector(83 downto 0);
             Y : in  std_logic_vector(83 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(83 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(52 downto 0);
signal YY_m6_c0 :  std_logic_vector(52 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c2 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c2, bh7_w0_0_c3, bh7_w0_0_c4 :  std_logic;
signal bh7_w1_0_c2, bh7_w1_0_c3, bh7_w1_0_c4 :  std_logic;
signal bh7_w2_0_c2, bh7_w2_0_c3, bh7_w2_0_c4 :  std_logic;
signal bh7_w3_0_c2, bh7_w3_0_c3, bh7_w3_0_c4 :  std_logic;
signal bh7_w4_0_c2, bh7_w4_0_c3, bh7_w4_0_c4 :  std_logic;
signal bh7_w5_0_c2, bh7_w5_0_c3, bh7_w5_0_c4 :  std_logic;
signal bh7_w6_0_c2, bh7_w6_0_c3, bh7_w6_0_c4 :  std_logic;
signal bh7_w7_0_c2, bh7_w7_0_c3, bh7_w7_0_c4 :  std_logic;
signal bh7_w8_0_c2, bh7_w8_0_c3, bh7_w8_0_c4 :  std_logic;
signal bh7_w9_0_c2, bh7_w9_0_c3, bh7_w9_0_c4 :  std_logic;
signal bh7_w10_0_c2, bh7_w10_0_c3, bh7_w10_0_c4 :  std_logic;
signal bh7_w11_0_c2, bh7_w11_0_c3, bh7_w11_0_c4 :  std_logic;
signal bh7_w12_0_c2, bh7_w12_0_c3, bh7_w12_0_c4 :  std_logic;
signal bh7_w13_0_c2, bh7_w13_0_c3, bh7_w13_0_c4 :  std_logic;
signal bh7_w14_0_c2, bh7_w14_0_c3, bh7_w14_0_c4 :  std_logic;
signal bh7_w15_0_c2, bh7_w15_0_c3, bh7_w15_0_c4 :  std_logic;
signal bh7_w16_0_c2, bh7_w16_0_c3, bh7_w16_0_c4 :  std_logic;
signal bh7_w17_0_c2 :  std_logic;
signal bh7_w18_0_c2 :  std_logic;
signal bh7_w19_0_c2 :  std_logic;
signal bh7_w20_0_c2 :  std_logic;
signal bh7_w21_0_c2 :  std_logic;
signal bh7_w22_0_c2 :  std_logic;
signal bh7_w23_0_c2 :  std_logic;
signal bh7_w24_0_c2 :  std_logic;
signal bh7_w25_0_c2 :  std_logic;
signal bh7_w26_0_c2 :  std_logic;
signal bh7_w27_0_c2 :  std_logic;
signal bh7_w28_0_c2 :  std_logic;
signal bh7_w29_0_c2 :  std_logic;
signal bh7_w30_0_c2 :  std_logic;
signal bh7_w31_0_c2 :  std_logic;
signal bh7_w32_0_c2 :  std_logic;
signal bh7_w33_0_c2 :  std_logic;
signal bh7_w34_0_c2 :  std_logic;
signal bh7_w35_0_c2 :  std_logic;
signal bh7_w36_0_c2 :  std_logic;
signal bh7_w37_0_c2 :  std_logic;
signal bh7_w38_0_c2 :  std_logic;
signal bh7_w39_0_c2 :  std_logic;
signal bh7_w40_0_c2 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(16 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_1_output_c2 :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w17_1_c2 :  std_logic;
signal bh7_w18_1_c2 :  std_logic;
signal bh7_w19_1_c2 :  std_logic;
signal bh7_w20_1_c2 :  std_logic;
signal bh7_w21_1_c2 :  std_logic;
signal bh7_w22_1_c2 :  std_logic;
signal bh7_w23_1_c2 :  std_logic;
signal bh7_w24_1_c2 :  std_logic;
signal bh7_w25_1_c2 :  std_logic;
signal bh7_w26_1_c2 :  std_logic;
signal bh7_w27_1_c2 :  std_logic;
signal bh7_w28_1_c2 :  std_logic;
signal bh7_w29_1_c2 :  std_logic;
signal bh7_w30_1_c2 :  std_logic;
signal bh7_w31_1_c2 :  std_logic;
signal bh7_w32_1_c2 :  std_logic;
signal bh7_w33_1_c2 :  std_logic;
signal bh7_w34_1_c2 :  std_logic;
signal bh7_w35_1_c2 :  std_logic;
signal bh7_w36_1_c2 :  std_logic;
signal bh7_w37_1_c2 :  std_logic;
signal bh7_w38_1_c2 :  std_logic;
signal bh7_w39_1_c2 :  std_logic;
signal bh7_w40_1_c2 :  std_logic;
signal bh7_w41_0_c2 :  std_logic;
signal bh7_w42_0_c2 :  std_logic;
signal bh7_w43_0_c2 :  std_logic;
signal bh7_w44_0_c2 :  std_logic;
signal bh7_w45_0_c2 :  std_logic;
signal bh7_w46_0_c2 :  std_logic;
signal bh7_w47_0_c2 :  std_logic;
signal bh7_w48_0_c2 :  std_logic;
signal bh7_w49_0_c2 :  std_logic;
signal bh7_w50_0_c2 :  std_logic;
signal bh7_w51_0_c2 :  std_logic;
signal bh7_w52_0_c2 :  std_logic;
signal bh7_w53_0_c2 :  std_logic;
signal bh7_w54_0_c2 :  std_logic;
signal bh7_w55_0_c2 :  std_logic;
signal bh7_w56_0_c2 :  std_logic;
signal bh7_w57_0_c2 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(16 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_2_output_c2 :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w34_2_c2 :  std_logic;
signal bh7_w35_2_c2 :  std_logic;
signal bh7_w36_2_c2 :  std_logic;
signal bh7_w37_2_c2 :  std_logic;
signal bh7_w38_2_c2 :  std_logic;
signal bh7_w39_2_c2 :  std_logic;
signal bh7_w40_2_c2 :  std_logic;
signal bh7_w41_1_c2 :  std_logic;
signal bh7_w42_1_c2 :  std_logic;
signal bh7_w43_1_c2 :  std_logic;
signal bh7_w44_1_c2 :  std_logic;
signal bh7_w45_1_c2 :  std_logic;
signal bh7_w46_1_c2 :  std_logic;
signal bh7_w47_1_c2 :  std_logic;
signal bh7_w48_1_c2 :  std_logic;
signal bh7_w49_1_c2 :  std_logic;
signal bh7_w50_1_c2 :  std_logic;
signal bh7_w51_1_c2 :  std_logic;
signal bh7_w52_1_c2 :  std_logic;
signal bh7_w53_1_c2 :  std_logic;
signal bh7_w54_1_c2 :  std_logic;
signal bh7_w55_1_c2 :  std_logic;
signal bh7_w56_1_c2 :  std_logic;
signal bh7_w57_1_c2 :  std_logic;
signal bh7_w58_0_c2 :  std_logic;
signal bh7_w59_0_c2, bh7_w59_0_c3 :  std_logic;
signal bh7_w60_0_c2, bh7_w60_0_c3 :  std_logic;
signal bh7_w61_0_c2, bh7_w61_0_c3 :  std_logic;
signal bh7_w62_0_c2, bh7_w62_0_c3 :  std_logic;
signal bh7_w63_0_c2 :  std_logic;
signal bh7_w64_0_c2, bh7_w64_0_c3 :  std_logic;
signal bh7_w65_0_c2, bh7_w65_0_c3 :  std_logic;
signal bh7_w66_0_c2 :  std_logic;
signal bh7_w67_0_c2, bh7_w67_0_c3 :  std_logic;
signal bh7_w68_0_c2 :  std_logic;
signal bh7_w69_0_c2, bh7_w69_0_c3 :  std_logic;
signal bh7_w70_0_c2, bh7_w70_0_c3 :  std_logic;
signal bh7_w71_0_c2 :  std_logic;
signal bh7_w72_0_c2, bh7_w72_0_c3 :  std_logic;
signal bh7_w73_0_c2 :  std_logic;
signal bh7_w74_0_c2, bh7_w74_0_c3 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w72_1_c0 :  std_logic;
signal bh7_w73_1_c0 :  std_logic;
signal bh7_w74_1_c0 :  std_logic;
signal bh7_w75_0_c0 :  std_logic;
signal bh7_w76_0_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_4_output_c0 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w69_1_c0 :  std_logic;
signal bh7_w70_1_c0 :  std_logic;
signal bh7_w71_1_c0 :  std_logic;
signal bh7_w72_2_c0 :  std_logic;
signal bh7_w73_2_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w66_1_c0 :  std_logic;
signal bh7_w67_1_c0 :  std_logic;
signal bh7_w68_1_c0 :  std_logic;
signal bh7_w69_2_c0 :  std_logic;
signal bh7_w70_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(1 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w63_1_c0 :  std_logic;
signal bh7_w64_1_c0 :  std_logic;
signal bh7_w65_1_c0 :  std_logic;
signal bh7_w66_2_c0 :  std_logic;
signal bh7_w67_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_7_output_c0 :  std_logic_vector(4 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_1_c0 :  std_logic;
signal bh7_w61_1_c0 :  std_logic;
signal bh7_w62_1_c0 :  std_logic;
signal bh7_w63_2_c0 :  std_logic;
signal bh7_w64_2_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(1 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_2_c0 :  std_logic;
signal bh7_w58_1_c0 :  std_logic;
signal bh7_w59_1_c0 :  std_logic;
signal bh7_w60_2_c0 :  std_logic;
signal bh7_w61_2_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(1 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_2_c0 :  std_logic;
signal bh7_w55_2_c0 :  std_logic;
signal bh7_w56_2_c0 :  std_logic;
signal bh7_w57_3_c0 :  std_logic;
signal bh7_w58_2_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_10_output_c0 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_2_c0 :  std_logic;
signal bh7_w52_2_c0 :  std_logic;
signal bh7_w53_2_c0 :  std_logic;
signal bh7_w54_3_c0 :  std_logic;
signal bh7_w55_3_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(16 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_11_output_c2 :  std_logic_vector(40 downto 0);
signal tile_11_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w24_2_c2 :  std_logic;
signal bh7_w25_2_c2, bh7_w25_2_c3 :  std_logic;
signal bh7_w26_2_c2 :  std_logic;
signal bh7_w27_2_c2, bh7_w27_2_c3 :  std_logic;
signal bh7_w28_2_c2 :  std_logic;
signal bh7_w29_2_c2, bh7_w29_2_c3 :  std_logic;
signal bh7_w30_2_c2 :  std_logic;
signal bh7_w31_2_c2, bh7_w31_2_c3 :  std_logic;
signal bh7_w32_2_c2 :  std_logic;
signal bh7_w33_2_c2, bh7_w33_2_c3 :  std_logic;
signal bh7_w34_3_c2 :  std_logic;
signal bh7_w35_3_c2 :  std_logic;
signal bh7_w36_3_c2 :  std_logic;
signal bh7_w37_3_c2 :  std_logic;
signal bh7_w38_3_c2 :  std_logic;
signal bh7_w39_3_c2 :  std_logic;
signal bh7_w40_3_c2 :  std_logic;
signal bh7_w41_2_c2 :  std_logic;
signal bh7_w42_2_c2 :  std_logic;
signal bh7_w43_2_c2 :  std_logic;
signal bh7_w44_2_c2 :  std_logic;
signal bh7_w45_2_c2 :  std_logic;
signal bh7_w46_2_c2 :  std_logic;
signal bh7_w47_2_c2 :  std_logic;
signal bh7_w48_2_c2 :  std_logic;
signal bh7_w49_2_c2 :  std_logic;
signal bh7_w50_2_c2 :  std_logic;
signal bh7_w51_3_c2 :  std_logic;
signal bh7_w52_3_c2 :  std_logic;
signal bh7_w53_3_c2 :  std_logic;
signal bh7_w54_4_c2 :  std_logic;
signal bh7_w55_4_c2 :  std_logic;
signal bh7_w56_3_c2 :  std_logic;
signal bh7_w57_4_c2 :  std_logic;
signal bh7_w58_3_c2 :  std_logic;
signal bh7_w59_2_c2, bh7_w59_2_c3 :  std_logic;
signal bh7_w60_3_c2, bh7_w60_3_c3 :  std_logic;
signal bh7_w61_3_c2, bh7_w61_3_c3 :  std_logic;
signal bh7_w62_2_c2, bh7_w62_2_c3 :  std_logic;
signal bh7_w63_3_c2 :  std_logic;
signal bh7_w64_3_c2, bh7_w64_3_c3 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(16 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_12_output_c2 :  std_logic_vector(40 downto 0);
signal tile_12_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w41_3_c2 :  std_logic;
signal bh7_w42_3_c2 :  std_logic;
signal bh7_w43_3_c2 :  std_logic;
signal bh7_w44_3_c2 :  std_logic;
signal bh7_w45_3_c2 :  std_logic;
signal bh7_w46_3_c2 :  std_logic;
signal bh7_w47_3_c2 :  std_logic;
signal bh7_w48_3_c2, bh7_w48_3_c3 :  std_logic;
signal bh7_w49_3_c2 :  std_logic;
signal bh7_w50_3_c2 :  std_logic;
signal bh7_w51_4_c2 :  std_logic;
signal bh7_w52_4_c2 :  std_logic;
signal bh7_w53_4_c2 :  std_logic;
signal bh7_w54_5_c2 :  std_logic;
signal bh7_w55_5_c2 :  std_logic;
signal bh7_w56_4_c2 :  std_logic;
signal bh7_w57_5_c2 :  std_logic;
signal bh7_w58_4_c2 :  std_logic;
signal bh7_w59_3_c2, bh7_w59_3_c3 :  std_logic;
signal bh7_w60_4_c2, bh7_w60_4_c3 :  std_logic;
signal bh7_w61_4_c2, bh7_w61_4_c3 :  std_logic;
signal bh7_w62_3_c2, bh7_w62_3_c3 :  std_logic;
signal bh7_w63_4_c2 :  std_logic;
signal bh7_w64_4_c2, bh7_w64_4_c3 :  std_logic;
signal bh7_w65_2_c2, bh7_w65_2_c3 :  std_logic;
signal bh7_w66_3_c2 :  std_logic;
signal bh7_w67_3_c2, bh7_w67_3_c3 :  std_logic;
signal bh7_w68_2_c2 :  std_logic;
signal bh7_w69_3_c2, bh7_w69_3_c3 :  std_logic;
signal bh7_w70_3_c2, bh7_w70_3_c3 :  std_logic;
signal bh7_w71_2_c2 :  std_logic;
signal bh7_w72_3_c2, bh7_w72_3_c3 :  std_logic;
signal bh7_w73_3_c2 :  std_logic;
signal bh7_w74_2_c2, bh7_w74_2_c3 :  std_logic;
signal bh7_w75_1_c2 :  std_logic;
signal bh7_w76_1_c2, bh7_w76_1_c3 :  std_logic;
signal bh7_w77_0_c2, bh7_w77_0_c3 :  std_logic;
signal bh7_w78_0_c2, bh7_w78_0_c3 :  std_logic;
signal bh7_w79_0_c2, bh7_w79_0_c3 :  std_logic;
signal bh7_w80_0_c2, bh7_w80_0_c3 :  std_logic;
signal bh7_w81_0_c2, bh7_w81_0_c3 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(16 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_13_output_c2 :  std_logic_vector(40 downto 0);
signal tile_13_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w58_5_c2, bh7_w58_5_c3 :  std_logic;
signal bh7_w59_4_c2, bh7_w59_4_c3 :  std_logic;
signal bh7_w60_5_c2, bh7_w60_5_c3 :  std_logic;
signal bh7_w61_5_c2, bh7_w61_5_c3 :  std_logic;
signal bh7_w62_4_c2, bh7_w62_4_c3 :  std_logic;
signal bh7_w63_5_c2, bh7_w63_5_c3 :  std_logic;
signal bh7_w64_5_c2, bh7_w64_5_c3 :  std_logic;
signal bh7_w65_3_c2, bh7_w65_3_c3 :  std_logic;
signal bh7_w66_4_c2 :  std_logic;
signal bh7_w67_4_c2, bh7_w67_4_c3 :  std_logic;
signal bh7_w68_3_c2 :  std_logic;
signal bh7_w69_4_c2, bh7_w69_4_c3 :  std_logic;
signal bh7_w70_4_c2, bh7_w70_4_c3 :  std_logic;
signal bh7_w71_3_c2 :  std_logic;
signal bh7_w72_4_c2, bh7_w72_4_c3 :  std_logic;
signal bh7_w73_4_c2 :  std_logic;
signal bh7_w74_3_c2, bh7_w74_3_c3 :  std_logic;
signal bh7_w75_2_c2, bh7_w75_2_c3 :  std_logic;
signal bh7_w76_2_c2, bh7_w76_2_c3 :  std_logic;
signal bh7_w77_1_c2, bh7_w77_1_c3 :  std_logic;
signal bh7_w78_1_c2, bh7_w78_1_c3 :  std_logic;
signal bh7_w79_1_c2, bh7_w79_1_c3 :  std_logic;
signal bh7_w80_1_c2, bh7_w80_1_c3 :  std_logic;
signal bh7_w81_1_c2, bh7_w81_1_c3 :  std_logic;
signal bh7_w82_0_c2, bh7_w82_0_c3 :  std_logic;
signal bh7_w83_0_c2, bh7_w83_0_c3 :  std_logic;
signal bh7_w84_0_c2, bh7_w84_0_c3 :  std_logic;
signal bh7_w85_0_c2, bh7_w85_0_c3 :  std_logic;
signal bh7_w86_0_c2, bh7_w86_0_c3 :  std_logic;
signal bh7_w87_0_c2, bh7_w87_0_c3 :  std_logic;
signal bh7_w88_0_c2, bh7_w88_0_c3 :  std_logic;
signal bh7_w89_0_c2, bh7_w89_0_c3 :  std_logic;
signal bh7_w90_0_c2, bh7_w90_0_c3 :  std_logic;
signal bh7_w91_0_c2, bh7_w91_0_c3 :  std_logic;
signal bh7_w92_0_c2, bh7_w92_0_c3 :  std_logic;
signal bh7_w93_0_c2, bh7_w93_0_c3 :  std_logic;
signal bh7_w94_0_c2, bh7_w94_0_c3 :  std_logic;
signal bh7_w95_0_c2, bh7_w95_0_c3 :  std_logic;
signal bh7_w96_0_c2, bh7_w96_0_c3 :  std_logic;
signal bh7_w97_0_c2, bh7_w97_0_c3 :  std_logic;
signal bh7_w98_0_c2, bh7_w98_0_c3 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(1 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_1_c0 :  std_logic;
signal bh7_w97_1_c0 :  std_logic;
signal bh7_w98_1_c0 :  std_logic;
signal bh7_w99_0_c0 :  std_logic;
signal bh7_w100_0_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_1_c0 :  std_logic;
signal bh7_w94_1_c0 :  std_logic;
signal bh7_w95_1_c0 :  std_logic;
signal bh7_w96_2_c0 :  std_logic;
signal bh7_w97_2_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_16_output_c0 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_1_c0 :  std_logic;
signal bh7_w91_1_c0 :  std_logic;
signal bh7_w92_1_c0 :  std_logic;
signal bh7_w93_2_c0 :  std_logic;
signal bh7_w94_2_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(1 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_1_c0 :  std_logic;
signal bh7_w88_1_c0 :  std_logic;
signal bh7_w89_1_c0 :  std_logic;
signal bh7_w90_2_c0 :  std_logic;
signal bh7_w91_2_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(1 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_1_c0 :  std_logic;
signal bh7_w85_1_c0 :  std_logic;
signal bh7_w86_1_c0 :  std_logic;
signal bh7_w87_2_c0 :  std_logic;
signal bh7_w88_2_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_19_output_c0 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w81_2_c0 :  std_logic;
signal bh7_w82_1_c0 :  std_logic;
signal bh7_w83_1_c0 :  std_logic;
signal bh7_w84_2_c0 :  std_logic;
signal bh7_w85_2_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(1 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w78_2_c0 :  std_logic;
signal bh7_w79_2_c0 :  std_logic;
signal bh7_w80_2_c0 :  std_logic;
signal bh7_w81_3_c0 :  std_logic;
signal bh7_w82_2_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(1 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w75_3_c0 :  std_logic;
signal bh7_w76_3_c0 :  std_logic;
signal bh7_w77_2_c0 :  std_logic;
signal bh7_w78_3_c0 :  std_logic;
signal bh7_w79_3_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_22_output_c0 :  std_logic_vector(0 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w68_4_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(3 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_23_output_c0 :  std_logic_vector(3 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w64_6_c0 :  std_logic;
signal bh7_w65_4_c0 :  std_logic;
signal bh7_w66_5_c0 :  std_logic;
signal bh7_w67_5_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(3 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_24_output_c0 :  std_logic_vector(3 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w60_6_c0 :  std_logic;
signal bh7_w61_6_c0 :  std_logic;
signal bh7_w62_5_c0 :  std_logic;
signal bh7_w63_6_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(3 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_25_output_c0 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w56_5_c0 :  std_logic;
signal bh7_w57_6_c0 :  std_logic;
signal bh7_w58_6_c0 :  std_logic;
signal bh7_w59_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(3 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_26_output_c0 :  std_logic_vector(3 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w52_5_c0 :  std_logic;
signal bh7_w53_5_c0 :  std_logic;
signal bh7_w54_6_c0 :  std_logic;
signal bh7_w55_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(1 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w65_5_c0 :  std_logic;
signal bh7_w66_6_c0 :  std_logic;
signal bh7_w67_6_c0 :  std_logic;
signal bh7_w68_5_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w62_6_c0 :  std_logic;
signal bh7_w63_7_c0 :  std_logic;
signal bh7_w64_7_c0 :  std_logic;
signal bh7_w65_6_c0 :  std_logic;
signal bh7_w66_7_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w59_6_c0 :  std_logic;
signal bh7_w60_7_c0 :  std_logic;
signal bh7_w61_7_c0 :  std_logic;
signal bh7_w62_7_c0 :  std_logic;
signal bh7_w63_8_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w56_6_c0 :  std_logic;
signal bh7_w57_7_c0 :  std_logic;
signal bh7_w58_7_c0 :  std_logic;
signal bh7_w59_7_c0 :  std_logic;
signal bh7_w60_8_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w53_6_c0 :  std_logic;
signal bh7_w54_7_c0 :  std_logic;
signal bh7_w55_7_c0 :  std_logic;
signal bh7_w56_7_c0 :  std_logic;
signal bh7_w57_8_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w50_4_c0 :  std_logic;
signal bh7_w51_5_c0 :  std_logic;
signal bh7_w52_6_c0 :  std_logic;
signal bh7_w53_7_c0 :  std_logic;
signal bh7_w54_8_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(1 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(3 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w63_9_c0 :  std_logic;
signal bh7_w64_8_c0 :  std_logic;
signal bh7_w65_7_c0 :  std_logic;
signal bh7_w66_8_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_9_c0 :  std_logic;
signal bh7_w61_8_c0 :  std_logic;
signal bh7_w62_8_c0, bh7_w62_8_c1 :  std_logic;
signal bh7_w63_10_c0 :  std_logic;
signal bh7_w64_9_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_9_c0 :  std_logic;
signal bh7_w58_8_c0 :  std_logic;
signal bh7_w59_8_c0, bh7_w59_8_c1 :  std_logic;
signal bh7_w60_10_c0 :  std_logic;
signal bh7_w61_9_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_9_c0 :  std_logic;
signal bh7_w55_8_c0 :  std_logic;
signal bh7_w56_8_c0, bh7_w56_8_c1 :  std_logic;
signal bh7_w57_10_c0 :  std_logic;
signal bh7_w58_9_c0 :  std_logic;
signal tile_37_X_c0 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_37_output_c0 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_6_c0 :  std_logic;
signal bh7_w52_7_c0 :  std_logic;
signal bh7_w53_8_c0 :  std_logic;
signal bh7_w54_10_c0 :  std_logic;
signal bh7_w55_9_c0 :  std_logic;
signal tile_38_X_c0 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_38_output_c0 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w48_4_c0, bh7_w48_4_c1, bh7_w48_4_c2 :  std_logic;
signal bh7_w49_4_c0 :  std_logic;
signal bh7_w50_5_c0 :  std_logic;
signal bh7_w51_7_c0 :  std_logic;
signal bh7_w52_8_c0 :  std_logic;
signal tile_39_X_c0 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_39_output_c0 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w85_3_c0 :  std_logic;
signal tile_40_X_c0 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_40_output_c0 :  std_logic_vector(3 downto 0);
signal tile_40_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w81_4_c0 :  std_logic;
signal bh7_w82_3_c0 :  std_logic;
signal bh7_w83_2_c0 :  std_logic;
signal bh7_w84_3_c0 :  std_logic;
signal tile_41_X_c0 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_41_output_c0 :  std_logic_vector(3 downto 0);
signal tile_41_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w77_3_c0 :  std_logic;
signal bh7_w78_4_c0 :  std_logic;
signal bh7_w79_4_c0 :  std_logic;
signal bh7_w80_3_c0 :  std_logic;
signal tile_42_X_c0 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_42_output_c0 :  std_logic_vector(3 downto 0);
signal tile_42_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w73_5_c0 :  std_logic;
signal bh7_w74_4_c0 :  std_logic;
signal bh7_w75_4_c0 :  std_logic;
signal bh7_w76_4_c0 :  std_logic;
signal tile_43_X_c0 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_43_output_c0 :  std_logic_vector(3 downto 0);
signal tile_43_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w69_5_c0 :  std_logic;
signal bh7_w70_5_c0 :  std_logic;
signal bh7_w71_4_c0 :  std_logic;
signal bh7_w72_5_c0 :  std_logic;
signal tile_44_X_c0 :  std_logic_vector(1 downto 0);
signal tile_44_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_44_output_c0 :  std_logic_vector(3 downto 0);
signal tile_44_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w82_4_c0 :  std_logic;
signal bh7_w83_3_c0 :  std_logic;
signal bh7_w84_4_c0 :  std_logic;
signal bh7_w85_4_c0 :  std_logic;
signal tile_45_X_c0 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_45_output_c0 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w79_5_c0 :  std_logic;
signal bh7_w80_4_c0 :  std_logic;
signal bh7_w81_5_c0 :  std_logic;
signal bh7_w82_5_c0 :  std_logic;
signal bh7_w83_4_c0 :  std_logic;
signal tile_46_X_c0 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_46_output_c0 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w76_5_c0 :  std_logic;
signal bh7_w77_4_c0 :  std_logic;
signal bh7_w78_5_c0 :  std_logic;
signal bh7_w79_6_c0 :  std_logic;
signal bh7_w80_5_c0 :  std_logic;
signal tile_47_X_c0 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_47_output_c0 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w73_6_c0 :  std_logic;
signal bh7_w74_5_c0 :  std_logic;
signal bh7_w75_5_c0 :  std_logic;
signal bh7_w76_6_c0 :  std_logic;
signal bh7_w77_5_c0 :  std_logic;
signal tile_48_X_c0 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_48_output_c0 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w70_6_c0 :  std_logic;
signal bh7_w71_5_c0 :  std_logic;
signal bh7_w72_6_c0 :  std_logic;
signal bh7_w73_7_c0 :  std_logic;
signal bh7_w74_6_c0 :  std_logic;
signal tile_49_X_c0 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_49_output_c0 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w67_7_c0 :  std_logic;
signal bh7_w68_6_c0 :  std_logic;
signal bh7_w69_6_c0 :  std_logic;
signal bh7_w70_7_c0 :  std_logic;
signal bh7_w71_6_c0 :  std_logic;
signal tile_50_X_c0 :  std_logic_vector(1 downto 0);
signal tile_50_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_50_output_c0 :  std_logic_vector(3 downto 0);
signal tile_50_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w80_6_c0 :  std_logic;
signal bh7_w81_6_c0 :  std_logic;
signal bh7_w82_6_c0 :  std_logic;
signal bh7_w83_5_c0 :  std_logic;
signal tile_51_X_c0 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_51_output_c0 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w77_6_c0 :  std_logic;
signal bh7_w78_6_c0 :  std_logic;
signal bh7_w79_7_c0 :  std_logic;
signal bh7_w80_7_c0 :  std_logic;
signal bh7_w81_7_c0 :  std_logic;
signal tile_52_X_c0 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_52_output_c0 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w74_7_c0 :  std_logic;
signal bh7_w75_6_c0 :  std_logic;
signal bh7_w76_7_c0 :  std_logic;
signal bh7_w77_7_c0 :  std_logic;
signal bh7_w78_7_c0 :  std_logic;
signal tile_53_X_c0 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_53_output_c0 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w71_7_c0 :  std_logic;
signal bh7_w72_7_c0 :  std_logic;
signal bh7_w73_8_c0 :  std_logic;
signal bh7_w74_8_c0 :  std_logic;
signal bh7_w75_7_c0 :  std_logic;
signal tile_54_X_c0 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_54_output_c0 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w68_7_c0 :  std_logic;
signal bh7_w69_7_c0 :  std_logic;
signal bh7_w70_8_c0 :  std_logic;
signal bh7_w71_8_c0 :  std_logic;
signal bh7_w72_8_c0 :  std_logic;
signal tile_55_X_c0 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_55_output_c0 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w65_8_c0 :  std_logic;
signal bh7_w66_9_c0, bh7_w66_9_c1 :  std_logic;
signal bh7_w67_8_c0 :  std_logic;
signal bh7_w68_8_c0 :  std_logic;
signal bh7_w69_8_c0 :  std_logic;
signal tile_56_X_c0 :  std_logic_vector(0 downto 0);
signal tile_56_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_56_output_c0 :  std_logic_vector(0 downto 0);
signal tile_56_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w102_0_c0 :  std_logic;
signal tile_57_X_c0 :  std_logic_vector(3 downto 0);
signal tile_57_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_57_output_c0 :  std_logic_vector(3 downto 0);
signal tile_57_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w98_2_c0 :  std_logic;
signal bh7_w99_1_c0 :  std_logic;
signal bh7_w100_1_c0 :  std_logic;
signal bh7_w101_0_c0 :  std_logic;
signal tile_58_X_c0 :  std_logic_vector(3 downto 0);
signal tile_58_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_58_output_c0 :  std_logic_vector(3 downto 0);
signal tile_58_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w94_3_c0 :  std_logic;
signal bh7_w95_2_c0 :  std_logic;
signal bh7_w96_3_c0 :  std_logic;
signal bh7_w97_3_c0 :  std_logic;
signal tile_59_X_c0 :  std_logic_vector(3 downto 0);
signal tile_59_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_59_output_c0 :  std_logic_vector(3 downto 0);
signal tile_59_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w90_3_c0 :  std_logic;
signal bh7_w91_3_c0 :  std_logic;
signal bh7_w92_2_c0 :  std_logic;
signal bh7_w93_3_c0 :  std_logic;
signal tile_60_X_c0 :  std_logic_vector(3 downto 0);
signal tile_60_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_60_output_c0 :  std_logic_vector(3 downto 0);
signal tile_60_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w86_2_c0 :  std_logic;
signal bh7_w87_3_c0 :  std_logic;
signal bh7_w88_3_c0 :  std_logic;
signal bh7_w89_2_c0 :  std_logic;
signal tile_61_X_c0 :  std_logic_vector(1 downto 0);
signal tile_61_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_61_output_c0 :  std_logic_vector(3 downto 0);
signal tile_61_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w99_2_c0 :  std_logic;
signal bh7_w100_2_c0 :  std_logic;
signal bh7_w101_1_c0 :  std_logic;
signal bh7_w102_1_c0 :  std_logic;
signal tile_62_X_c0 :  std_logic_vector(2 downto 0);
signal tile_62_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_62_output_c0 :  std_logic_vector(4 downto 0);
signal tile_62_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_4_c0 :  std_logic;
signal bh7_w97_4_c0 :  std_logic;
signal bh7_w98_3_c0 :  std_logic;
signal bh7_w99_3_c0 :  std_logic;
signal bh7_w100_3_c0 :  std_logic;
signal tile_63_X_c0 :  std_logic_vector(2 downto 0);
signal tile_63_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_63_output_c0 :  std_logic_vector(4 downto 0);
signal tile_63_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_4_c0 :  std_logic;
signal bh7_w94_4_c0 :  std_logic;
signal bh7_w95_3_c0 :  std_logic;
signal bh7_w96_5_c0 :  std_logic;
signal bh7_w97_5_c0 :  std_logic;
signal tile_64_X_c0 :  std_logic_vector(2 downto 0);
signal tile_64_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_64_output_c0 :  std_logic_vector(4 downto 0);
signal tile_64_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_4_c0 :  std_logic;
signal bh7_w91_4_c0 :  std_logic;
signal bh7_w92_3_c0 :  std_logic;
signal bh7_w93_5_c0 :  std_logic;
signal bh7_w94_5_c0 :  std_logic;
signal tile_65_X_c0 :  std_logic_vector(2 downto 0);
signal tile_65_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_65_output_c0 :  std_logic_vector(4 downto 0);
signal tile_65_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_4_c0 :  std_logic;
signal bh7_w88_4_c0 :  std_logic;
signal bh7_w89_3_c0 :  std_logic;
signal bh7_w90_5_c0 :  std_logic;
signal bh7_w91_5_c0 :  std_logic;
signal tile_66_X_c0 :  std_logic_vector(2 downto 0);
signal tile_66_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_66_output_c0 :  std_logic_vector(4 downto 0);
signal tile_66_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_5_c0 :  std_logic;
signal bh7_w85_5_c0 :  std_logic;
signal bh7_w86_3_c0 :  std_logic;
signal bh7_w87_5_c0 :  std_logic;
signal bh7_w88_5_c0 :  std_logic;
signal tile_67_X_c0 :  std_logic_vector(1 downto 0);
signal tile_67_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_67_output_c0 :  std_logic_vector(3 downto 0);
signal tile_67_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w97_6_c0 :  std_logic;
signal bh7_w98_4_c0 :  std_logic;
signal bh7_w99_4_c0 :  std_logic;
signal bh7_w100_4_c0 :  std_logic;
signal tile_68_X_c0 :  std_logic_vector(2 downto 0);
signal tile_68_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_68_output_c0 :  std_logic_vector(4 downto 0);
signal tile_68_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w94_6_c0 :  std_logic;
signal bh7_w95_4_c0 :  std_logic;
signal bh7_w96_6_c0 :  std_logic;
signal bh7_w97_7_c0, bh7_w97_7_c1 :  std_logic;
signal bh7_w98_5_c0 :  std_logic;
signal tile_69_X_c0 :  std_logic_vector(2 downto 0);
signal tile_69_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_69_output_c0 :  std_logic_vector(4 downto 0);
signal tile_69_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w91_6_c0 :  std_logic;
signal bh7_w92_4_c0 :  std_logic;
signal bh7_w93_6_c0 :  std_logic;
signal bh7_w94_7_c0, bh7_w94_7_c1 :  std_logic;
signal bh7_w95_5_c0 :  std_logic;
signal tile_70_X_c0 :  std_logic_vector(2 downto 0);
signal tile_70_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_70_output_c0 :  std_logic_vector(4 downto 0);
signal tile_70_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w88_6_c0 :  std_logic;
signal bh7_w89_4_c0 :  std_logic;
signal bh7_w90_6_c0 :  std_logic;
signal bh7_w91_7_c0, bh7_w91_7_c1 :  std_logic;
signal bh7_w92_5_c0 :  std_logic;
signal tile_71_X_c0 :  std_logic_vector(2 downto 0);
signal tile_71_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_71_output_c0 :  std_logic_vector(4 downto 0);
signal tile_71_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w85_6_c0 :  std_logic;
signal bh7_w86_4_c0 :  std_logic;
signal bh7_w87_6_c0 :  std_logic;
signal bh7_w88_7_c0, bh7_w88_7_c1 :  std_logic;
signal bh7_w89_5_c0 :  std_logic;
signal tile_72_X_c0 :  std_logic_vector(2 downto 0);
signal tile_72_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_72_output_c0 :  std_logic_vector(4 downto 0);
signal tile_72_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w82_7_c0, bh7_w82_7_c1 :  std_logic;
signal bh7_w83_6_c0 :  std_logic;
signal bh7_w84_6_c0 :  std_logic;
signal bh7_w85_7_c0, bh7_w85_7_c1 :  std_logic;
signal bh7_w86_5_c0 :  std_logic;
signal tile_73_X_c0 :  std_logic_vector(1 downto 0);
signal tile_73_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_73_output_c0 :  std_logic_vector(3 downto 0);
signal tile_73_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w102_2_c0 :  std_logic;
signal bh7_w103_0_c0 :  std_logic;
signal bh7_w104_0_c0, bh7_w104_0_c1 :  std_logic;
signal bh7_w105_0_c0, bh7_w105_0_c1 :  std_logic;
signal tile_74_X_c0 :  std_logic_vector(1 downto 0);
signal tile_74_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_74_output_c0 :  std_logic_vector(4 downto 0);
signal tile_74_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w99_5_c0 :  std_logic;
signal bh7_w100_5_c0 :  std_logic;
signal bh7_w101_2_c0 :  std_logic;
signal bh7_w102_3_c0 :  std_logic;
signal bh7_w103_1_c0, bh7_w103_1_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid323_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid323_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w49_5_c1 :  std_logic;
signal bh7_w50_6_c1 :  std_logic;
signal bh7_w51_8_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c0, Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid327_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid327_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_9_c1 :  std_logic;
signal bh7_w52_9_c1 :  std_logic;
signal bh7_w53_9_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c0, Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid329_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid329_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_10_c1 :  std_logic;
signal bh7_w53_10_c1 :  std_logic;
signal bh7_w54_11_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c0, Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid331_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid331_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_11_c1 :  std_logic;
signal bh7_w54_12_c1 :  std_logic;
signal bh7_w55_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c0, Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid335_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_13_c1 :  std_logic;
signal bh7_w55_11_c1 :  std_logic;
signal bh7_w56_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c0, Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid337_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_12_c1 :  std_logic;
signal bh7_w56_10_c1 :  std_logic;
signal bh7_w57_11_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c0, Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid339_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid339_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_11_c1 :  std_logic;
signal bh7_w57_12_c1 :  std_logic;
signal bh7_w58_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c0, Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid341_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_13_c1 :  std_logic;
signal bh7_w58_11_c1 :  std_logic;
signal bh7_w59_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c0, Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid343_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_12_c1 :  std_logic;
signal bh7_w59_10_c1 :  std_logic;
signal bh7_w60_11_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c0, Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid345_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid345_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_11_c1 :  std_logic;
signal bh7_w60_12_c1 :  std_logic;
signal bh7_w61_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c0, Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid347_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_13_c1 :  std_logic;
signal bh7_w61_11_c1 :  std_logic;
signal bh7_w62_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c0, Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid349_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w61_12_c1 :  std_logic;
signal bh7_w62_10_c1 :  std_logic;
signal bh7_w63_11_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c0, Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid351_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid351_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_11_c1 :  std_logic;
signal bh7_w63_12_c1 :  std_logic;
signal bh7_w64_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c0, Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid353_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w63_13_c1 :  std_logic;
signal bh7_w64_11_c1 :  std_logic;
signal bh7_w65_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c0, Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid355_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_12_c1 :  std_logic;
signal bh7_w65_10_c1 :  std_logic;
signal bh7_w66_10_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c0, Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid357_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_11_c1 :  std_logic;
signal bh7_w66_11_c1 :  std_logic;
signal bh7_w67_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c0, Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid359_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_12_c1 :  std_logic;
signal bh7_w67_10_c1 :  std_logic;
signal bh7_w68_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c0, Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid361_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_11_c1 :  std_logic;
signal bh7_w68_10_c1 :  std_logic;
signal bh7_w69_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c0, Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid363_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_11_c1 :  std_logic;
signal bh7_w69_10_c1 :  std_logic;
signal bh7_w70_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c0, Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid365_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w69_11_c1 :  std_logic;
signal bh7_w70_10_c1 :  std_logic;
signal bh7_w71_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c0, Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid367_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_11_c1 :  std_logic;
signal bh7_w71_10_c1 :  std_logic;
signal bh7_w72_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c0, Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid369_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w71_11_c1 :  std_logic;
signal bh7_w72_10_c1 :  std_logic;
signal bh7_w73_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c0, Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid371_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_11_c1 :  std_logic;
signal bh7_w73_10_c1 :  std_logic;
signal bh7_w74_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c0, Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid373_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w73_11_c1 :  std_logic;
signal bh7_w74_10_c1 :  std_logic;
signal bh7_w75_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c0, Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid375_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_11_c1 :  std_logic;
signal bh7_w75_9_c1 :  std_logic;
signal bh7_w76_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c0, Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid377_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w75_10_c1 :  std_logic;
signal bh7_w76_9_c1 :  std_logic;
signal bh7_w77_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c0, Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid379_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_10_c1 :  std_logic;
signal bh7_w77_9_c1 :  std_logic;
signal bh7_w78_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c0, Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid381_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w77_10_c1 :  std_logic;
signal bh7_w78_9_c1 :  std_logic;
signal bh7_w79_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c0, Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid383_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_10_c1 :  std_logic;
signal bh7_w79_9_c1 :  std_logic;
signal bh7_w80_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c0, Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid385_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w79_10_c1 :  std_logic;
signal bh7_w80_9_c1 :  std_logic;
signal bh7_w81_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c0, Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid387_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_10_c1 :  std_logic;
signal bh7_w81_9_c1 :  std_logic;
signal bh7_w82_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c0, Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid389_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w81_10_c1 :  std_logic;
signal bh7_w82_9_c1 :  std_logic;
signal bh7_w83_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c0, Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid391_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_10_c1 :  std_logic;
signal bh7_w83_8_c1 :  std_logic;
signal bh7_w84_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c0, Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid393_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w83_9_c1 :  std_logic;
signal bh7_w84_8_c1 :  std_logic;
signal bh7_w85_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c0, Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid395_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_9_c1 :  std_logic;
signal bh7_w85_9_c1 :  std_logic;
signal bh7_w86_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c0, Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid397_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w85_10_c1 :  std_logic;
signal bh7_w86_7_c1 :  std_logic;
signal bh7_w87_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c0, Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid401_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_8_c1 :  std_logic;
signal bh7_w87_8_c1 :  std_logic;
signal bh7_w88_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c0, Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid403_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w87_9_c1 :  std_logic;
signal bh7_w88_9_c1 :  std_logic;
signal bh7_w89_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c0, Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid405_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_10_c1 :  std_logic;
signal bh7_w89_7_c1 :  std_logic;
signal bh7_w90_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c0, Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid407_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w89_8_c1 :  std_logic;
signal bh7_w90_8_c1 :  std_logic;
signal bh7_w91_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c0, Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid409_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_9_c1 :  std_logic;
signal bh7_w91_9_c1 :  std_logic;
signal bh7_w92_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c0, Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid411_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_10_c1 :  std_logic;
signal bh7_w92_7_c1 :  std_logic;
signal bh7_w93_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c0, Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid413_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_8_c1 :  std_logic;
signal bh7_w93_8_c1 :  std_logic;
signal bh7_w94_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c0, Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid415_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w93_9_c1 :  std_logic;
signal bh7_w94_9_c1 :  std_logic;
signal bh7_w95_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c0, Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid417_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_10_c1 :  std_logic;
signal bh7_w95_7_c1 :  std_logic;
signal bh7_w96_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c0, Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid419_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w95_8_c1 :  std_logic;
signal bh7_w96_8_c1 :  std_logic;
signal bh7_w97_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c0, Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid421_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w96_9_c1 :  std_logic;
signal bh7_w97_9_c1 :  std_logic;
signal bh7_w98_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c0, Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid423_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_10_c1 :  std_logic;
signal bh7_w98_7_c1 :  std_logic;
signal bh7_w99_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c0, Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid425_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_8_c1 :  std_logic;
signal bh7_w99_7_c1 :  std_logic;
signal bh7_w100_6_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c0, Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid427_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w99_8_c1 :  std_logic;
signal bh7_w100_7_c1 :  std_logic;
signal bh7_w101_3_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c0, Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid429_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_8_c1 :  std_logic;
signal bh7_w101_4_c1 :  std_logic;
signal bh7_w102_4_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c0, Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid433_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w101_5_c1 :  std_logic;
signal bh7_w102_5_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c0, Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid435_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid435_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w102_6_c1 :  std_logic;
signal bh7_w103_2_c1 :  std_logic;
signal bh7_w104_1_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c0, Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid437_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid437_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_10_c1 :  std_logic;
signal bh7_w52_11_c1 :  std_logic;
signal bh7_w53_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_copy438_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid439_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid439_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_13_c1 :  std_logic;
signal bh7_w54_14_c1 :  std_logic;
signal bh7_w55_13_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_copy440_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid441_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w55_14_c1 :  std_logic;
signal bh7_w56_12_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_copy442_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid443_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_13_c1 :  std_logic;
signal bh7_w57_14_c1 :  std_logic;
signal bh7_w58_13_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_copy444_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid445_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w57_15_c1 :  std_logic;
signal bh7_w58_14_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_copy446_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid447_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w58_15_c1 :  std_logic;
signal bh7_w59_12_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_copy448_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid449_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_13_c1 :  std_logic;
signal bh7_w60_14_c1 :  std_logic;
signal bh7_w61_13_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_copy450_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid451_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w60_15_c1 :  std_logic;
signal bh7_w61_14_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_copy452_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid453_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w61_15_c1 :  std_logic;
signal bh7_w62_12_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_copy454_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid455_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_13_c1 :  std_logic;
signal bh7_w63_14_c1 :  std_logic;
signal bh7_w64_13_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_copy456_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid457_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w63_15_c1 :  std_logic;
signal bh7_w64_14_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_copy458_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid459_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid459_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_15_c1 :  std_logic;
signal bh7_w65_12_c1 :  std_logic;
signal bh7_w66_13_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_copy460_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid461_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_14_c1 :  std_logic;
signal bh7_w67_12_c1 :  std_logic;
signal bh7_w68_12_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_copy462_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid463_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w67_13_c1 :  std_logic;
signal bh7_w68_13_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_copy464_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid465_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid465_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_14_c1 :  std_logic;
signal bh7_w69_12_c1 :  std_logic;
signal bh7_w70_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_copy466_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid467_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid467_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_13_c1 :  std_logic;
signal bh7_w71_12_c1 :  std_logic;
signal bh7_w72_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_copy468_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid469_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid469_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_13_c1 :  std_logic;
signal bh7_w73_12_c1 :  std_logic;
signal bh7_w74_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_copy470_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid471_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid471_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_13_c1 :  std_logic;
signal bh7_w75_11_c1 :  std_logic;
signal bh7_w76_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_copy472_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid473_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid473_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_12_c1 :  std_logic;
signal bh7_w77_11_c1 :  std_logic;
signal bh7_w78_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_copy474_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid475_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid475_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_12_c1 :  std_logic;
signal bh7_w79_11_c1 :  std_logic;
signal bh7_w80_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_copy476_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid477_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid477_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_12_c1 :  std_logic;
signal bh7_w81_11_c1 :  std_logic;
signal bh7_w82_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_copy478_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid479_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_12_c1 :  std_logic;
signal bh7_w83_10_c1 :  std_logic;
signal bh7_w84_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_copy480_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid481_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w83_11_c1 :  std_logic;
signal bh7_w84_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_copy482_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid483_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w84_12_c1 :  std_logic;
signal bh7_w85_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_copy484_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid485_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w85_12_c1 :  std_logic;
signal bh7_w86_9_c1 :  std_logic;
signal bh7_w87_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_copy486_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid487_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w86_10_c1 :  std_logic;
signal bh7_w87_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_copy488_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid489_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w87_12_c1 :  std_logic;
signal bh7_w88_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_copy490_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid491_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_12_c1 :  std_logic;
signal bh7_w89_9_c1 :  std_logic;
signal bh7_w90_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_copy492_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid493_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w89_10_c1 :  std_logic;
signal bh7_w90_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_copy494_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid495_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w90_12_c1 :  std_logic;
signal bh7_w91_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_copy496_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid497_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_12_c1 :  std_logic;
signal bh7_w92_9_c1 :  std_logic;
signal bh7_w93_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_copy498_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid499_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w92_10_c1 :  std_logic;
signal bh7_w93_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_copy500_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid501_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w93_12_c1 :  std_logic;
signal bh7_w94_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_copy502_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid503_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_12_c1 :  std_logic;
signal bh7_w95_9_c1 :  std_logic;
signal bh7_w96_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_copy504_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid505_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w95_10_c1 :  std_logic;
signal bh7_w96_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_copy506_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid507_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w96_12_c1 :  std_logic;
signal bh7_w97_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_copy508_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid509_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_12_c1 :  std_logic;
signal bh7_w98_9_c1 :  std_logic;
signal bh7_w99_9_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_copy510_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid511_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w98_10_c1 :  std_logic;
signal bh7_w99_10_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_copy512_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid513_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid513_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w99_11_c1 :  std_logic;
signal bh7_w100_9_c1 :  std_logic;
signal bh7_w101_6_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_copy514_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid515_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid515_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w101_7_c1 :  std_logic;
signal bh7_w102_7_c1 :  std_logic;
signal bh7_w103_3_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_copy516_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid517_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid517_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_4_c1 :  std_logic;
signal bh7_w104_2_c1 :  std_logic;
signal bh7_w105_1_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_copy518_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid519_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid519_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w53_14_c2 :  std_logic;
signal bh7_w54_15_c2 :  std_logic;
signal bh7_w55_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c1, Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid521_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid521_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w55_16_c2 :  std_logic;
signal bh7_w56_14_c2 :  std_logic;
signal bh7_w57_16_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c1, Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid523_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w57_17_c2 :  std_logic;
signal bh7_w58_16_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c1, Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid525_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid525_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w58_17_c2 :  std_logic;
signal bh7_w59_14_c2 :  std_logic;
signal bh7_w60_16_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c1, Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid527_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w60_17_c2 :  std_logic;
signal bh7_w61_16_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c1, Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid529_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid529_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w61_17_c2 :  std_logic;
signal bh7_w62_14_c2 :  std_logic;
signal bh7_w63_16_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c1, Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid531_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w63_17_c2 :  std_logic;
signal bh7_w64_16_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c1, Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid533_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid533_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w64_17_c2 :  std_logic;
signal bh7_w65_13_c2 :  std_logic;
signal bh7_w66_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c1, Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid535_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid535_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w66_16_c2 :  std_logic;
signal bh7_w67_14_c2 :  std_logic;
signal bh7_w68_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c1, Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid537_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid537_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w68_16_c2 :  std_logic;
signal bh7_w69_13_c2 :  std_logic;
signal bh7_w70_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c1, Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid539_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid539_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w70_15_c2 :  std_logic;
signal bh7_w71_13_c2 :  std_logic;
signal bh7_w72_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c1, Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid541_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid541_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w72_15_c2 :  std_logic;
signal bh7_w73_13_c2 :  std_logic;
signal bh7_w74_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c1, Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid543_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid543_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w74_15_c2 :  std_logic;
signal bh7_w75_12_c2 :  std_logic;
signal bh7_w76_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c1, Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid545_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid545_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w76_14_c2 :  std_logic;
signal bh7_w77_12_c2 :  std_logic;
signal bh7_w78_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c1, Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid547_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid547_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w78_14_c2 :  std_logic;
signal bh7_w79_12_c2 :  std_logic;
signal bh7_w80_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c1, Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid549_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid549_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w80_14_c2 :  std_logic;
signal bh7_w81_12_c2 :  std_logic;
signal bh7_w82_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c1, Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid551_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid551_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w82_14_c2 :  std_logic;
signal bh7_w83_12_c2 :  std_logic;
signal bh7_w84_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c1, Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid553_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid553_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w84_14_c2 :  std_logic;
signal bh7_w85_13_c2 :  std_logic;
signal bh7_w86_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c1, Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid555_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w86_12_c2 :  std_logic;
signal bh7_w87_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c1, Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid557_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid557_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w87_14_c2 :  std_logic;
signal bh7_w88_13_c2 :  std_logic;
signal bh7_w89_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c1, Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid559_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w89_12_c2 :  std_logic;
signal bh7_w90_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c1, Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid561_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid561_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w90_14_c2 :  std_logic;
signal bh7_w91_13_c2 :  std_logic;
signal bh7_w92_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c1, Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid563_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w92_12_c2 :  std_logic;
signal bh7_w93_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c1, Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid565_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid565_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w93_14_c2 :  std_logic;
signal bh7_w94_13_c2 :  std_logic;
signal bh7_w95_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c1, Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid567_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w95_12_c2 :  std_logic;
signal bh7_w96_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c1, Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid569_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid569_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w96_14_c2 :  std_logic;
signal bh7_w97_13_c2 :  std_logic;
signal bh7_w98_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c1, Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid571_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w98_12_c2 :  std_logic;
signal bh7_w99_12_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c1, Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid573_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid573_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w99_13_c2 :  std_logic;
signal bh7_w100_10_c2 :  std_logic;
signal bh7_w101_8_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c1, Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid575_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid575_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w101_9_c2 :  std_logic;
signal bh7_w102_8_c2 :  std_logic;
signal bh7_w103_5_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c1, Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid577_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid577_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w103_6_c2 :  std_logic;
signal bh7_w104_3_c2 :  std_logic;
signal bh7_w105_2_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c1, Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid579_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w105_3_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c1, Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c2 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid581_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid581_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w55_17_c2 :  std_logic;
signal bh7_w56_15_c2 :  std_logic;
signal bh7_w57_18_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_copy582_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid583_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid583_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w57_19_c2 :  std_logic;
signal bh7_w58_18_c2 :  std_logic;
signal bh7_w59_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_copy584_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid585_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid585_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w60_18_c2 :  std_logic;
signal bh7_w61_18_c2, bh7_w61_18_c3 :  std_logic;
signal bh7_w62_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_copy586_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid587_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid587_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w63_18_c2 :  std_logic;
signal bh7_w64_18_c2, bh7_w64_18_c3 :  std_logic;
signal bh7_w65_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_copy588_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid589_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid589_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w66_17_c2 :  std_logic;
signal bh7_w67_15_c2, bh7_w67_15_c3 :  std_logic;
signal bh7_w68_17_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_copy590_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid591_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid591_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w68_18_c2 :  std_logic;
signal bh7_w69_14_c2 :  std_logic;
signal bh7_w70_16_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_copy592_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid593_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid593_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w70_17_c2 :  std_logic;
signal bh7_w71_14_c2 :  std_logic;
signal bh7_w72_16_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_copy594_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid595_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid595_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w72_17_c2 :  std_logic;
signal bh7_w73_14_c2 :  std_logic;
signal bh7_w74_16_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_copy596_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid597_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid597_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w74_17_c2 :  std_logic;
signal bh7_w75_13_c2 :  std_logic;
signal bh7_w76_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_copy598_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid599_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid599_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w76_16_c2 :  std_logic;
signal bh7_w77_13_c2 :  std_logic;
signal bh7_w78_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_copy600_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid601_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid601_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w78_16_c2 :  std_logic;
signal bh7_w79_13_c2 :  std_logic;
signal bh7_w80_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_copy602_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid603_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid603_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w80_16_c2 :  std_logic;
signal bh7_w81_13_c2 :  std_logic;
signal bh7_w82_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_copy604_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid605_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid605_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w82_16_c2 :  std_logic;
signal bh7_w83_13_c2 :  std_logic;
signal bh7_w84_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_copy606_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid607_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid607_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w84_16_c2 :  std_logic;
signal bh7_w85_14_c2 :  std_logic;
signal bh7_w86_13_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_copy608_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid609_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid609_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w86_14_c2 :  std_logic;
signal bh7_w87_15_c2 :  std_logic;
signal bh7_w88_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_copy610_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid611_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid611_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w89_13_c2 :  std_logic;
signal bh7_w90_15_c2, bh7_w90_15_c3 :  std_logic;
signal bh7_w91_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_copy612_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid613_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid613_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w92_13_c2 :  std_logic;
signal bh7_w93_15_c2, bh7_w93_15_c3 :  std_logic;
signal bh7_w94_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_copy614_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid615_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid615_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w95_13_c2 :  std_logic;
signal bh7_w96_15_c2, bh7_w96_15_c3 :  std_logic;
signal bh7_w97_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_copy616_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid617_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid617_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w98_13_c2 :  std_logic;
signal bh7_w99_14_c2, bh7_w99_14_c3 :  std_logic;
signal bh7_w100_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_copy618_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid619_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid619_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w101_10_c2 :  std_logic;
signal bh7_w102_9_c2, bh7_w102_9_c3 :  std_logic;
signal bh7_w103_7_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_copy620_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid621_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid621_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w103_8_c2 :  std_logic;
signal bh7_w104_4_c2 :  std_logic;
signal bh7_w105_4_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_copy622_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid623_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w105_5_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_copy624_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid625_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid625_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w57_20_c3 :  std_logic;
signal bh7_w58_19_c3 :  std_logic;
signal bh7_w59_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c2, Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid627_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid627_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w59_17_c3 :  std_logic;
signal bh7_w60_19_c3 :  std_logic;
signal bh7_w61_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c2, Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid629_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid629_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w62_16_c3 :  std_logic;
signal bh7_w63_19_c3 :  std_logic;
signal bh7_w64_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c2, Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid631_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid631_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w65_15_c3 :  std_logic;
signal bh7_w66_18_c3 :  std_logic;
signal bh7_w67_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c2, Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid633_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid633_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w68_19_c3 :  std_logic;
signal bh7_w69_15_c3 :  std_logic;
signal bh7_w70_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c2, Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid635_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid635_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w70_19_c3 :  std_logic;
signal bh7_w71_15_c3 :  std_logic;
signal bh7_w72_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c2, Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid637_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid637_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w72_19_c3 :  std_logic;
signal bh7_w73_15_c3 :  std_logic;
signal bh7_w74_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c2, Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid639_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid639_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w74_19_c3 :  std_logic;
signal bh7_w75_14_c3 :  std_logic;
signal bh7_w76_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c2, Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid641_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid641_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w76_18_c3 :  std_logic;
signal bh7_w77_14_c3 :  std_logic;
signal bh7_w78_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c2, Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid643_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid643_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w78_18_c3 :  std_logic;
signal bh7_w79_14_c3 :  std_logic;
signal bh7_w80_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c2, Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid645_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid645_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w80_18_c3 :  std_logic;
signal bh7_w81_14_c3 :  std_logic;
signal bh7_w82_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c2, Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid647_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid647_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w82_18_c3 :  std_logic;
signal bh7_w83_14_c3 :  std_logic;
signal bh7_w84_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c2, Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid649_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid649_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w84_18_c3 :  std_logic;
signal bh7_w85_15_c3 :  std_logic;
signal bh7_w86_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c2, Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid651_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid651_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w86_16_c3 :  std_logic;
signal bh7_w87_16_c3 :  std_logic;
signal bh7_w88_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c2, Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid653_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid653_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w88_16_c3 :  std_logic;
signal bh7_w89_14_c3 :  std_logic;
signal bh7_w90_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c2, Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid655_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid655_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w91_15_c3 :  std_logic;
signal bh7_w92_14_c3 :  std_logic;
signal bh7_w93_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c2, Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid657_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid657_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w94_15_c3 :  std_logic;
signal bh7_w95_14_c3 :  std_logic;
signal bh7_w96_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c2, Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid659_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid659_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w97_15_c3 :  std_logic;
signal bh7_w98_14_c3 :  std_logic;
signal bh7_w99_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c2, Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid661_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid661_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w100_12_c3 :  std_logic;
signal bh7_w101_11_c3 :  std_logic;
signal bh7_w102_10_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c2, Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid663_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid663_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w103_9_c3 :  std_logic;
signal bh7_w104_5_c3 :  std_logic;
signal bh7_w105_6_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c2, Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid665_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w105_7_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c2, Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid667_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid667_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c3, bh7_w17_2_c4 :  std_logic;
signal bh7_w18_2_c3, bh7_w18_2_c4 :  std_logic;
signal bh7_w19_2_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c2, Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid669_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid669_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w19_3_c3 :  std_logic;
signal bh7_w20_2_c3 :  std_logic;
signal bh7_w21_2_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c2, Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid671_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid671_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w21_3_c3 :  std_logic;
signal bh7_w22_2_c3 :  std_logic;
signal bh7_w23_2_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c2, Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid673_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w23_3_c3 :  std_logic;
signal bh7_w24_3_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c2, Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid675_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid675_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w24_4_c3 :  std_logic;
signal bh7_w25_3_c3 :  std_logic;
signal bh7_w26_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c2, Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid677_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid677_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w26_4_c3 :  std_logic;
signal bh7_w27_3_c3 :  std_logic;
signal bh7_w28_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c2, Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid679_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid679_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w28_4_c3 :  std_logic;
signal bh7_w29_3_c3 :  std_logic;
signal bh7_w30_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c2, Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid681_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid681_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w30_4_c3 :  std_logic;
signal bh7_w31_3_c3 :  std_logic;
signal bh7_w32_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c2, Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid683_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid683_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w32_4_c3 :  std_logic;
signal bh7_w33_3_c3 :  std_logic;
signal bh7_w34_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c2, Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid685_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid685_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w34_5_c3 :  std_logic;
signal bh7_w35_4_c3 :  std_logic;
signal bh7_w36_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c2, Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid687_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w35_5_c3 :  std_logic;
signal bh7_w36_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c2, Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid689_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid689_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w36_6_c3 :  std_logic;
signal bh7_w37_4_c3 :  std_logic;
signal bh7_w38_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c2, Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid691_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w37_5_c3 :  std_logic;
signal bh7_w38_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c2, Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid693_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid693_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w38_6_c3 :  std_logic;
signal bh7_w39_4_c3 :  std_logic;
signal bh7_w40_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c2, Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid695_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w39_5_c3 :  std_logic;
signal bh7_w40_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c2, Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid697_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid697_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w40_6_c3 :  std_logic;
signal bh7_w41_4_c3 :  std_logic;
signal bh7_w42_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c2, Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid699_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w41_5_c3 :  std_logic;
signal bh7_w42_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c2, Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid701_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid701_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w42_6_c3 :  std_logic;
signal bh7_w43_4_c3 :  std_logic;
signal bh7_w44_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c2, Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid703_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w43_5_c3 :  std_logic;
signal bh7_w44_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c2, Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid705_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid705_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w44_6_c3 :  std_logic;
signal bh7_w45_4_c3 :  std_logic;
signal bh7_w46_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c2, Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid707_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w45_5_c3 :  std_logic;
signal bh7_w46_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c2, Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid709_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid709_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w46_6_c3 :  std_logic;
signal bh7_w47_4_c3 :  std_logic;
signal bh7_w48_5_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c2, Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid711_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w47_5_c3 :  std_logic;
signal bh7_w48_6_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c2, Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid713_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w48_7_c3 :  std_logic;
signal bh7_w49_6_c3 :  std_logic;
signal bh7_w50_7_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c2, Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid715_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w49_7_c3 :  std_logic;
signal bh7_w50_8_c3 :  std_logic;
signal bh7_w51_11_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c2, Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid717_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w50_9_c3 :  std_logic;
signal bh7_w51_12_c3 :  std_logic;
signal bh7_w52_12_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c2, Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid719_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w51_13_c3 :  std_logic;
signal bh7_w52_13_c3 :  std_logic;
signal bh7_w53_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c2, Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid721_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid721_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w52_14_c3 :  std_logic;
signal bh7_w53_16_c3 :  std_logic;
signal bh7_w54_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c2, Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid723_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid723_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w53_17_c3 :  std_logic;
signal bh7_w54_17_c3 :  std_logic;
signal bh7_w55_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c2, Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid725_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid725_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w54_18_c3 :  std_logic;
signal bh7_w55_19_c3 :  std_logic;
signal bh7_w56_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c2, Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid727_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid727_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w55_20_c3 :  std_logic;
signal bh7_w56_17_c3 :  std_logic;
signal bh7_w57_21_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c2, Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c2, Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid729_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w56_18_c3 :  std_logic;
signal bh7_w57_22_c3 :  std_logic;
signal bh7_w58_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_copy730_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c2, Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid731_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w57_23_c3, bh7_w57_23_c4 :  std_logic;
signal bh7_w58_21_c3 :  std_logic;
signal bh7_w59_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_copy732_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid733_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w58_22_c3 :  std_logic;
signal bh7_w59_19_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c2, Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c3 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid735_In0_c3 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w59_20_c3 :  std_logic;
signal bh7_w60_20_c3 :  std_logic;
signal bh7_w61_20_c3 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_copy736_c3 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid737_In0_c3 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w60_21_c3 :  std_logic;
signal bh7_w61_21_c3 :  std_logic;
signal bh7_w62_17_c3 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_copy738_c3 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid739_In0_c3 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w61_22_c3 :  std_logic;
signal bh7_w62_18_c3 :  std_logic;
signal bh7_w63_20_c3 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_copy740_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid741_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid741_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w62_19_c3 :  std_logic;
signal bh7_w63_21_c3 :  std_logic;
signal bh7_w64_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_copy742_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid743_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w63_22_c3 :  std_logic;
signal bh7_w64_21_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c2, Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c3 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid745_In0_c3 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w64_22_c3 :  std_logic;
signal bh7_w65_16_c3 :  std_logic;
signal bh7_w66_19_c3 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_copy746_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid747_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid747_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w65_17_c3 :  std_logic;
signal bh7_w66_20_c3 :  std_logic;
signal bh7_w67_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_copy748_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid749_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w66_21_c3 :  std_logic;
signal bh7_w67_18_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c2, Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid751_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid751_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w67_19_c3 :  std_logic;
signal bh7_w68_20_c3 :  std_logic;
signal bh7_w69_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_copy752_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid753_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w68_21_c3, bh7_w68_21_c4 :  std_logic;
signal bh7_w69_17_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c2, Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid755_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid755_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w69_18_c3 :  std_logic;
signal bh7_w70_20_c3 :  std_logic;
signal bh7_w71_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_copy756_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid757_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid757_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w70_21_c3 :  std_logic;
signal bh7_w71_17_c3 :  std_logic;
signal bh7_w72_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_copy758_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid759_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w71_18_c3 :  std_logic;
signal bh7_w72_21_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c2, Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid761_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid761_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w72_22_c3 :  std_logic;
signal bh7_w73_16_c3 :  std_logic;
signal bh7_w74_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_copy762_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid763_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w73_17_c3, bh7_w73_17_c4 :  std_logic;
signal bh7_w74_21_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c2, Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid765_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w74_22_c3 :  std_logic;
signal bh7_w75_15_c3 :  std_logic;
signal bh7_w76_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_copy766_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid767_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid767_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w74_23_c3 :  std_logic;
signal bh7_w75_16_c3, bh7_w75_16_c4 :  std_logic;
signal bh7_w76_20_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_copy768_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid769_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w76_21_c3 :  std_logic;
signal bh7_w77_15_c3 :  std_logic;
signal bh7_w78_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_copy770_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid771_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w77_16_c3 :  std_logic;
signal bh7_w78_20_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_copy772_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid773_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w78_21_c3 :  std_logic;
signal bh7_w79_15_c3 :  std_logic;
signal bh7_w80_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_copy774_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid775_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w79_16_c3 :  std_logic;
signal bh7_w80_20_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_copy776_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid777_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w80_21_c3 :  std_logic;
signal bh7_w81_15_c3 :  std_logic;
signal bh7_w82_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_copy778_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid779_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w81_16_c3 :  std_logic;
signal bh7_w82_20_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_copy780_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid781_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid781_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w82_21_c3 :  std_logic;
signal bh7_w83_15_c3, bh7_w83_15_c4 :  std_logic;
signal bh7_w84_19_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_copy782_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid783_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid783_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w84_20_c3 :  std_logic;
signal bh7_w85_16_c3 :  std_logic;
signal bh7_w86_17_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_copy784_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid785_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid785_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w86_18_c3 :  std_logic;
signal bh7_w87_17_c3 :  std_logic;
signal bh7_w88_17_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_copy786_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid787_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid787_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w88_18_c3 :  std_logic;
signal bh7_w89_15_c3 :  std_logic;
signal bh7_w90_17_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_copy788_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid789_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid789_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w90_18_c3 :  std_logic;
signal bh7_w91_16_c3 :  std_logic;
signal bh7_w92_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_copy790_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid791_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w92_16_c3 :  std_logic;
signal bh7_w93_17_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_copy792_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid793_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid793_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w93_18_c3 :  std_logic;
signal bh7_w94_16_c3, bh7_w94_16_c4 :  std_logic;
signal bh7_w95_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_copy794_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid795_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w95_16_c3 :  std_logic;
signal bh7_w96_17_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_copy796_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid797_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid797_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w96_18_c3 :  std_logic;
signal bh7_w97_16_c3, bh7_w97_16_c4 :  std_logic;
signal bh7_w98_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_copy798_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid799_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid799_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w98_16_c3 :  std_logic;
signal bh7_w99_16_c3 :  std_logic;
signal bh7_w100_13_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_copy800_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid801_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid801_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w102_11_c3, bh7_w102_11_c4 :  std_logic;
signal bh7_w103_10_c3 :  std_logic;
signal bh7_w104_6_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_copy802_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid803_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w105_8_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_copy804_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid805_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid805_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w19_4_c3, bh7_w19_4_c4 :  std_logic;
signal bh7_w20_3_c3, bh7_w20_3_c4 :  std_logic;
signal bh7_w21_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_copy806_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid807_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid807_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w21_5_c3 :  std_logic;
signal bh7_w22_3_c3 :  std_logic;
signal bh7_w23_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_copy808_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid809_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid809_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w23_5_c3 :  std_logic;
signal bh7_w24_5_c3 :  std_logic;
signal bh7_w25_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_copy810_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid811_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid811_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w25_5_c3 :  std_logic;
signal bh7_w26_5_c3 :  std_logic;
signal bh7_w27_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_copy812_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid813_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid813_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w27_5_c3 :  std_logic;
signal bh7_w28_5_c3 :  std_logic;
signal bh7_w29_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_copy814_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid815_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid815_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w29_5_c3 :  std_logic;
signal bh7_w30_5_c3 :  std_logic;
signal bh7_w31_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_copy816_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid817_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid817_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w31_5_c3 :  std_logic;
signal bh7_w32_5_c3 :  std_logic;
signal bh7_w33_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_copy818_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid819_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid819_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w33_5_c3 :  std_logic;
signal bh7_w34_6_c3 :  std_logic;
signal bh7_w35_6_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_copy820_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid821_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w35_7_c3 :  std_logic;
signal bh7_w36_7_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_copy822_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid823_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid823_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w36_8_c3 :  std_logic;
signal bh7_w37_6_c3, bh7_w37_6_c4 :  std_logic;
signal bh7_w38_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_copy824_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid825_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid825_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w38_8_c3 :  std_logic;
signal bh7_w39_6_c3 :  std_logic;
signal bh7_w40_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_copy826_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid827_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid827_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w40_8_c3 :  std_logic;
signal bh7_w41_6_c3 :  std_logic;
signal bh7_w42_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_copy828_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid829_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid829_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w42_8_c3 :  std_logic;
signal bh7_w43_6_c3 :  std_logic;
signal bh7_w44_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_copy830_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid831_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid831_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w44_8_c3 :  std_logic;
signal bh7_w45_6_c3 :  std_logic;
signal bh7_w46_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_copy832_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid833_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid833_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w46_8_c3 :  std_logic;
signal bh7_w47_6_c3 :  std_logic;
signal bh7_w48_8_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_copy834_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid835_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid835_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w48_9_c3 :  std_logic;
signal bh7_w49_8_c3 :  std_logic;
signal bh7_w50_10_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_copy836_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid837_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid837_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w50_11_c3 :  std_logic;
signal bh7_w51_14_c3 :  std_logic;
signal bh7_w52_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_copy838_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid839_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid839_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w52_16_c3 :  std_logic;
signal bh7_w53_18_c3 :  std_logic;
signal bh7_w54_19_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_copy840_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid841_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid841_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w54_20_c3 :  std_logic;
signal bh7_w55_21_c3 :  std_logic;
signal bh7_w56_19_c3, bh7_w56_19_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_copy842_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid843_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid843_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w56_20_c4 :  std_logic;
signal bh7_w57_24_c4 :  std_logic;
signal bh7_w58_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c3, Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid845_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w58_24_c4 :  std_logic;
signal bh7_w59_21_c4 :  std_logic;
signal bh7_w60_22_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c3, Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid847_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid847_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w59_22_c4 :  std_logic;
signal bh7_w60_23_c4 :  std_logic;
signal bh7_w61_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c3, Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid849_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w61_24_c4 :  std_logic;
signal bh7_w62_20_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c3, Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid851_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid851_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w62_21_c4 :  std_logic;
signal bh7_w63_23_c4 :  std_logic;
signal bh7_w64_23_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c3, Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid853_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c0, Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c1, Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c2, Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w63_24_c4 :  std_logic;
signal bh7_w64_24_c4 :  std_logic;
signal bh7_w65_18_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c3, Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid855_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid855_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w64_25_c4 :  std_logic;
signal bh7_w65_19_c4 :  std_logic;
signal bh7_w66_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c3, Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid857_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w66_23_c4 :  std_logic;
signal bh7_w67_20_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c3, Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid859_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid859_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w67_21_c4 :  std_logic;
signal bh7_w68_22_c4 :  std_logic;
signal bh7_w69_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c3, Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid861_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid861_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w69_20_c4 :  std_logic;
signal bh7_w70_22_c4 :  std_logic;
signal bh7_w71_19_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c3, Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid863_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w71_20_c4 :  std_logic;
signal bh7_w72_23_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c3, Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid865_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid865_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w72_24_c4 :  std_logic;
signal bh7_w73_18_c4 :  std_logic;
signal bh7_w74_24_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c3, Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid867_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid867_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w74_25_c4 :  std_logic;
signal bh7_w75_17_c4 :  std_logic;
signal bh7_w76_22_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c3, Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid869_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid869_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w76_23_c4 :  std_logic;
signal bh7_w77_17_c4 :  std_logic;
signal bh7_w78_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c3, Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid871_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid871_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w78_23_c4 :  std_logic;
signal bh7_w79_17_c4 :  std_logic;
signal bh7_w80_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c3, Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid873_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid873_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w80_23_c4 :  std_logic;
signal bh7_w81_17_c4 :  std_logic;
signal bh7_w82_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c3, Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid875_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w82_23_c4 :  std_logic;
signal bh7_w83_16_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c3, Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid877_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid877_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w84_21_c4 :  std_logic;
signal bh7_w85_17_c4 :  std_logic;
signal bh7_w86_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c3, Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid879_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid879_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w86_20_c4 :  std_logic;
signal bh7_w87_18_c4 :  std_logic;
signal bh7_w88_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c3, Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid881_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid881_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w88_20_c4 :  std_logic;
signal bh7_w89_16_c4 :  std_logic;
signal bh7_w90_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c3, Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid883_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid883_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w90_20_c4 :  std_logic;
signal bh7_w91_17_c4 :  std_logic;
signal bh7_w92_17_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c3, Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid885_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid885_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w92_18_c4 :  std_logic;
signal bh7_w93_19_c4 :  std_logic;
signal bh7_w94_17_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c3, Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid887_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid887_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w95_17_c4 :  std_logic;
signal bh7_w96_19_c4 :  std_logic;
signal bh7_w97_17_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c3, Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid889_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid889_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w98_17_c4 :  std_logic;
signal bh7_w99_17_c4 :  std_logic;
signal bh7_w100_14_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c3, Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid891_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid891_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w100_15_c4 :  std_logic;
signal bh7_w101_12_c4 :  std_logic;
signal bh7_w102_12_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c3, Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid893_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid893_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w104_7_c4 :  std_logic;
signal bh7_w105_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c3, Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid895_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid895_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c4 :  std_logic;
signal bh7_w22_4_c4 :  std_logic;
signal bh7_w23_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c3, Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid897_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid897_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w23_7_c4 :  std_logic;
signal bh7_w24_6_c4 :  std_logic;
signal bh7_w25_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c3, Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid899_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid899_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w25_7_c4 :  std_logic;
signal bh7_w26_6_c4 :  std_logic;
signal bh7_w27_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c3, Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid901_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid901_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w27_7_c4 :  std_logic;
signal bh7_w28_6_c4 :  std_logic;
signal bh7_w29_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c3, Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid903_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid903_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w29_7_c4 :  std_logic;
signal bh7_w30_6_c4 :  std_logic;
signal bh7_w31_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c3, Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid905_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid905_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w31_7_c4 :  std_logic;
signal bh7_w32_6_c4 :  std_logic;
signal bh7_w33_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c3, Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid907_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid907_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w33_7_c4 :  std_logic;
signal bh7_w34_7_c4 :  std_logic;
signal bh7_w35_8_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c3, Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid909_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid909_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c4 :  std_logic;
signal bh7_w36_9_c4 :  std_logic;
signal bh7_w37_7_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c3, Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid911_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid911_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c4 :  std_logic;
signal bh7_w39_7_c4 :  std_logic;
signal bh7_w40_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c3, Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid913_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid913_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w40_10_c4 :  std_logic;
signal bh7_w41_7_c4 :  std_logic;
signal bh7_w42_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c3, Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid915_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid915_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w42_10_c4 :  std_logic;
signal bh7_w43_7_c4 :  std_logic;
signal bh7_w44_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c3, Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid917_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid917_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w44_10_c4 :  std_logic;
signal bh7_w45_7_c4 :  std_logic;
signal bh7_w46_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c3, Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid919_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid919_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w46_10_c4 :  std_logic;
signal bh7_w47_7_c4 :  std_logic;
signal bh7_w48_10_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c3, Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid921_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid921_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w48_11_c4 :  std_logic;
signal bh7_w49_9_c4 :  std_logic;
signal bh7_w50_12_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c3, Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid923_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid923_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w50_13_c4 :  std_logic;
signal bh7_w51_15_c4 :  std_logic;
signal bh7_w52_17_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c3, Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid925_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid925_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w52_18_c4 :  std_logic;
signal bh7_w53_19_c4 :  std_logic;
signal bh7_w54_21_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c3, Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid927_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid927_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w54_22_c4 :  std_logic;
signal bh7_w55_22_c4 :  std_logic;
signal bh7_w56_21_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c3, Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid929_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid929_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w56_22_c4 :  std_logic;
signal bh7_w57_25_c4 :  std_logic;
signal bh7_w58_25_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_copy930_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid931_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid931_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w58_26_c4 :  std_logic;
signal bh7_w59_23_c4 :  std_logic;
signal bh7_w60_24_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_copy932_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid933_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid933_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w60_25_c4 :  std_logic;
signal bh7_w61_25_c4 :  std_logic;
signal bh7_w62_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_copy934_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid935_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid935_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w62_23_c4 :  std_logic;
signal bh7_w63_25_c4 :  std_logic;
signal bh7_w64_26_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_copy936_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid937_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid937_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w64_27_c4 :  std_logic;
signal bh7_w65_20_c4 :  std_logic;
signal bh7_w66_24_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_copy938_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid939_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid939_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w66_25_c4 :  std_logic;
signal bh7_w67_22_c4 :  std_logic;
signal bh7_w68_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_copy940_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid941_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid941_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w68_24_c4 :  std_logic;
signal bh7_w69_21_c4 :  std_logic;
signal bh7_w70_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_copy942_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid943_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid943_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w71_21_c4 :  std_logic;
signal bh7_w72_25_c4 :  std_logic;
signal bh7_w73_19_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_copy944_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid945_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid945_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w73_20_c4 :  std_logic;
signal bh7_w74_26_c4 :  std_logic;
signal bh7_w75_18_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_copy946_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid947_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid947_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w75_19_c4 :  std_logic;
signal bh7_w76_24_c4 :  std_logic;
signal bh7_w77_18_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_copy948_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid949_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid949_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w78_24_c4 :  std_logic;
signal bh7_w79_18_c4 :  std_logic;
signal bh7_w80_24_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_copy950_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid951_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid951_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w80_25_c4 :  std_logic;
signal bh7_w81_18_c4 :  std_logic;
signal bh7_w82_24_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_copy952_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid953_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid953_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w82_25_c4 :  std_logic;
signal bh7_w83_17_c4 :  std_logic;
signal bh7_w84_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_copy954_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid955_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid955_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w86_21_c4 :  std_logic;
signal bh7_w87_19_c4 :  std_logic;
signal bh7_w88_21_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_copy956_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid957_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid957_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w88_22_c4 :  std_logic;
signal bh7_w89_17_c4 :  std_logic;
signal bh7_w90_21_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_copy958_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid959_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid959_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w90_22_c4 :  std_logic;
signal bh7_w91_18_c4 :  std_logic;
signal bh7_w92_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_copy960_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid961_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid961_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w92_20_c4 :  std_logic;
signal bh7_w93_20_c4 :  std_logic;
signal bh7_w94_18_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_copy962_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid963_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid963_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w94_19_c4 :  std_logic;
signal bh7_w95_18_c4 :  std_logic;
signal bh7_w96_20_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_copy964_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid965_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid965_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w97_18_c4 :  std_logic;
signal bh7_w98_18_c4 :  std_logic;
signal bh7_w99_18_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_copy966_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid967_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid967_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w100_16_c4 :  std_logic;
signal bh7_w101_13_c4 :  std_logic;
signal bh7_w102_13_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_copy968_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid969_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c3, Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w102_14_c4 :  std_logic;
signal bh7_w103_11_c4 :  std_logic;
signal bh7_w104_8_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_copy970_c4 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_22_c4, tmp_bitheapResult_bh7_22_c5, tmp_bitheapResult_bh7_22_c6, tmp_bitheapResult_bh7_22_c7, tmp_bitheapResult_bh7_22_c8, tmp_bitheapResult_bh7_22_c9, tmp_bitheapResult_bh7_22_c10, tmp_bitheapResult_bh7_22_c11, tmp_bitheapResult_bh7_22_c12, tmp_bitheapResult_bh7_22_c13, tmp_bitheapResult_bh7_22_c14, tmp_bitheapResult_bh7_22_c15, tmp_bitheapResult_bh7_22_c16, tmp_bitheapResult_bh7_22_c17, tmp_bitheapResult_bh7_22_c18, tmp_bitheapResult_bh7_22_c19, tmp_bitheapResult_bh7_22_c20, tmp_bitheapResult_bh7_22_c21, tmp_bitheapResult_bh7_22_c22, tmp_bitheapResult_bh7_22_c23, tmp_bitheapResult_bh7_22_c24, tmp_bitheapResult_bh7_22_c25, tmp_bitheapResult_bh7_22_c26, tmp_bitheapResult_bh7_22_c27, tmp_bitheapResult_bh7_22_c28, tmp_bitheapResult_bh7_22_c29, tmp_bitheapResult_bh7_22_c30, tmp_bitheapResult_bh7_22_c31, tmp_bitheapResult_bh7_22_c32, tmp_bitheapResult_bh7_22_c33 :  std_logic_vector(22 downto 0);
signal bitheapFinalAdd_bh7_In0_c4 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_In1_c4 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c33 :  std_logic_vector(83 downto 0);
signal bitheapResult_bh7_c33 :  std_logic_vector(105 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w62_8_c1 <= bh7_w62_8_c0;
               bh7_w59_8_c1 <= bh7_w59_8_c0;
               bh7_w56_8_c1 <= bh7_w56_8_c0;
               bh7_w48_4_c1 <= bh7_w48_4_c0;
               bh7_w66_9_c1 <= bh7_w66_9_c0;
               bh7_w97_7_c1 <= bh7_w97_7_c0;
               bh7_w94_7_c1 <= bh7_w94_7_c0;
               bh7_w91_7_c1 <= bh7_w91_7_c0;
               bh7_w88_7_c1 <= bh7_w88_7_c0;
               bh7_w82_7_c1 <= bh7_w82_7_c0;
               bh7_w85_7_c1 <= bh7_w85_7_c0;
               bh7_w104_0_c1 <= bh7_w104_0_c0;
               bh7_w105_0_c1 <= bh7_w105_0_c0;
               bh7_w103_1_c1 <= bh7_w103_1_c0;
               Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c0;
               Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c0;
               Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c0;
            end if;
            if ce_2 = '1' then
               bh7_w48_4_c2 <= bh7_w48_4_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c1;
            end if;
            if ce_3 = '1' then
               bh7_w0_0_c3 <= bh7_w0_0_c2;
               bh7_w1_0_c3 <= bh7_w1_0_c2;
               bh7_w2_0_c3 <= bh7_w2_0_c2;
               bh7_w3_0_c3 <= bh7_w3_0_c2;
               bh7_w4_0_c3 <= bh7_w4_0_c2;
               bh7_w5_0_c3 <= bh7_w5_0_c2;
               bh7_w6_0_c3 <= bh7_w6_0_c2;
               bh7_w7_0_c3 <= bh7_w7_0_c2;
               bh7_w8_0_c3 <= bh7_w8_0_c2;
               bh7_w9_0_c3 <= bh7_w9_0_c2;
               bh7_w10_0_c3 <= bh7_w10_0_c2;
               bh7_w11_0_c3 <= bh7_w11_0_c2;
               bh7_w12_0_c3 <= bh7_w12_0_c2;
               bh7_w13_0_c3 <= bh7_w13_0_c2;
               bh7_w14_0_c3 <= bh7_w14_0_c2;
               bh7_w15_0_c3 <= bh7_w15_0_c2;
               bh7_w16_0_c3 <= bh7_w16_0_c2;
               bh7_w59_0_c3 <= bh7_w59_0_c2;
               bh7_w60_0_c3 <= bh7_w60_0_c2;
               bh7_w61_0_c3 <= bh7_w61_0_c2;
               bh7_w62_0_c3 <= bh7_w62_0_c2;
               bh7_w64_0_c3 <= bh7_w64_0_c2;
               bh7_w65_0_c3 <= bh7_w65_0_c2;
               bh7_w67_0_c3 <= bh7_w67_0_c2;
               bh7_w69_0_c3 <= bh7_w69_0_c2;
               bh7_w70_0_c3 <= bh7_w70_0_c2;
               bh7_w72_0_c3 <= bh7_w72_0_c2;
               bh7_w74_0_c3 <= bh7_w74_0_c2;
               bh7_w25_2_c3 <= bh7_w25_2_c2;
               bh7_w27_2_c3 <= bh7_w27_2_c2;
               bh7_w29_2_c3 <= bh7_w29_2_c2;
               bh7_w31_2_c3 <= bh7_w31_2_c2;
               bh7_w33_2_c3 <= bh7_w33_2_c2;
               bh7_w59_2_c3 <= bh7_w59_2_c2;
               bh7_w60_3_c3 <= bh7_w60_3_c2;
               bh7_w61_3_c3 <= bh7_w61_3_c2;
               bh7_w62_2_c3 <= bh7_w62_2_c2;
               bh7_w64_3_c3 <= bh7_w64_3_c2;
               bh7_w48_3_c3 <= bh7_w48_3_c2;
               bh7_w59_3_c3 <= bh7_w59_3_c2;
               bh7_w60_4_c3 <= bh7_w60_4_c2;
               bh7_w61_4_c3 <= bh7_w61_4_c2;
               bh7_w62_3_c3 <= bh7_w62_3_c2;
               bh7_w64_4_c3 <= bh7_w64_4_c2;
               bh7_w65_2_c3 <= bh7_w65_2_c2;
               bh7_w67_3_c3 <= bh7_w67_3_c2;
               bh7_w69_3_c3 <= bh7_w69_3_c2;
               bh7_w70_3_c3 <= bh7_w70_3_c2;
               bh7_w72_3_c3 <= bh7_w72_3_c2;
               bh7_w74_2_c3 <= bh7_w74_2_c2;
               bh7_w76_1_c3 <= bh7_w76_1_c2;
               bh7_w77_0_c3 <= bh7_w77_0_c2;
               bh7_w78_0_c3 <= bh7_w78_0_c2;
               bh7_w79_0_c3 <= bh7_w79_0_c2;
               bh7_w80_0_c3 <= bh7_w80_0_c2;
               bh7_w81_0_c3 <= bh7_w81_0_c2;
               bh7_w58_5_c3 <= bh7_w58_5_c2;
               bh7_w59_4_c3 <= bh7_w59_4_c2;
               bh7_w60_5_c3 <= bh7_w60_5_c2;
               bh7_w61_5_c3 <= bh7_w61_5_c2;
               bh7_w62_4_c3 <= bh7_w62_4_c2;
               bh7_w63_5_c3 <= bh7_w63_5_c2;
               bh7_w64_5_c3 <= bh7_w64_5_c2;
               bh7_w65_3_c3 <= bh7_w65_3_c2;
               bh7_w67_4_c3 <= bh7_w67_4_c2;
               bh7_w69_4_c3 <= bh7_w69_4_c2;
               bh7_w70_4_c3 <= bh7_w70_4_c2;
               bh7_w72_4_c3 <= bh7_w72_4_c2;
               bh7_w74_3_c3 <= bh7_w74_3_c2;
               bh7_w75_2_c3 <= bh7_w75_2_c2;
               bh7_w76_2_c3 <= bh7_w76_2_c2;
               bh7_w77_1_c3 <= bh7_w77_1_c2;
               bh7_w78_1_c3 <= bh7_w78_1_c2;
               bh7_w79_1_c3 <= bh7_w79_1_c2;
               bh7_w80_1_c3 <= bh7_w80_1_c2;
               bh7_w81_1_c3 <= bh7_w81_1_c2;
               bh7_w82_0_c3 <= bh7_w82_0_c2;
               bh7_w83_0_c3 <= bh7_w83_0_c2;
               bh7_w84_0_c3 <= bh7_w84_0_c2;
               bh7_w85_0_c3 <= bh7_w85_0_c2;
               bh7_w86_0_c3 <= bh7_w86_0_c2;
               bh7_w87_0_c3 <= bh7_w87_0_c2;
               bh7_w88_0_c3 <= bh7_w88_0_c2;
               bh7_w89_0_c3 <= bh7_w89_0_c2;
               bh7_w90_0_c3 <= bh7_w90_0_c2;
               bh7_w91_0_c3 <= bh7_w91_0_c2;
               bh7_w92_0_c3 <= bh7_w92_0_c2;
               bh7_w93_0_c3 <= bh7_w93_0_c2;
               bh7_w94_0_c3 <= bh7_w94_0_c2;
               bh7_w95_0_c3 <= bh7_w95_0_c2;
               bh7_w96_0_c3 <= bh7_w96_0_c2;
               bh7_w97_0_c3 <= bh7_w97_0_c2;
               bh7_w98_0_c3 <= bh7_w98_0_c2;
               bh7_w61_18_c3 <= bh7_w61_18_c2;
               bh7_w64_18_c3 <= bh7_w64_18_c2;
               bh7_w67_15_c3 <= bh7_w67_15_c2;
               bh7_w90_15_c3 <= bh7_w90_15_c2;
               bh7_w93_15_c3 <= bh7_w93_15_c2;
               bh7_w96_15_c3 <= bh7_w96_15_c2;
               bh7_w99_14_c3 <= bh7_w99_14_c2;
               bh7_w102_9_c3 <= bh7_w102_9_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c2;
            end if;
            if ce_4 = '1' then
               bh7_w0_0_c4 <= bh7_w0_0_c3;
               bh7_w1_0_c4 <= bh7_w1_0_c3;
               bh7_w2_0_c4 <= bh7_w2_0_c3;
               bh7_w3_0_c4 <= bh7_w3_0_c3;
               bh7_w4_0_c4 <= bh7_w4_0_c3;
               bh7_w5_0_c4 <= bh7_w5_0_c3;
               bh7_w6_0_c4 <= bh7_w6_0_c3;
               bh7_w7_0_c4 <= bh7_w7_0_c3;
               bh7_w8_0_c4 <= bh7_w8_0_c3;
               bh7_w9_0_c4 <= bh7_w9_0_c3;
               bh7_w10_0_c4 <= bh7_w10_0_c3;
               bh7_w11_0_c4 <= bh7_w11_0_c3;
               bh7_w12_0_c4 <= bh7_w12_0_c3;
               bh7_w13_0_c4 <= bh7_w13_0_c3;
               bh7_w14_0_c4 <= bh7_w14_0_c3;
               bh7_w15_0_c4 <= bh7_w15_0_c3;
               bh7_w16_0_c4 <= bh7_w16_0_c3;
               bh7_w17_2_c4 <= bh7_w17_2_c3;
               bh7_w18_2_c4 <= bh7_w18_2_c3;
               bh7_w57_23_c4 <= bh7_w57_23_c3;
               bh7_w68_21_c4 <= bh7_w68_21_c3;
               bh7_w73_17_c4 <= bh7_w73_17_c3;
               bh7_w75_16_c4 <= bh7_w75_16_c3;
               bh7_w83_15_c4 <= bh7_w83_15_c3;
               bh7_w94_16_c4 <= bh7_w94_16_c3;
               bh7_w97_16_c4 <= bh7_w97_16_c3;
               bh7_w102_11_c4 <= bh7_w102_11_c3;
               bh7_w19_4_c4 <= bh7_w19_4_c3;
               bh7_w20_3_c4 <= bh7_w20_3_c3;
               bh7_w37_6_c4 <= bh7_w37_6_c3;
               bh7_w56_19_c4 <= bh7_w56_19_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c3;
            end if;
            if ce_5 = '1' then
               tmp_bitheapResult_bh7_22_c5 <= tmp_bitheapResult_bh7_22_c4;
            end if;
            if ce_6 = '1' then
               tmp_bitheapResult_bh7_22_c6 <= tmp_bitheapResult_bh7_22_c5;
            end if;
            if ce_7 = '1' then
               tmp_bitheapResult_bh7_22_c7 <= tmp_bitheapResult_bh7_22_c6;
            end if;
            if ce_8 = '1' then
               tmp_bitheapResult_bh7_22_c8 <= tmp_bitheapResult_bh7_22_c7;
            end if;
            if ce_9 = '1' then
               tmp_bitheapResult_bh7_22_c9 <= tmp_bitheapResult_bh7_22_c8;
            end if;
            if ce_10 = '1' then
               tmp_bitheapResult_bh7_22_c10 <= tmp_bitheapResult_bh7_22_c9;
            end if;
            if ce_11 = '1' then
               tmp_bitheapResult_bh7_22_c11 <= tmp_bitheapResult_bh7_22_c10;
            end if;
            if ce_12 = '1' then
               tmp_bitheapResult_bh7_22_c12 <= tmp_bitheapResult_bh7_22_c11;
            end if;
            if ce_13 = '1' then
               tmp_bitheapResult_bh7_22_c13 <= tmp_bitheapResult_bh7_22_c12;
            end if;
            if ce_14 = '1' then
               tmp_bitheapResult_bh7_22_c14 <= tmp_bitheapResult_bh7_22_c13;
            end if;
            if ce_15 = '1' then
               tmp_bitheapResult_bh7_22_c15 <= tmp_bitheapResult_bh7_22_c14;
            end if;
            if ce_16 = '1' then
               tmp_bitheapResult_bh7_22_c16 <= tmp_bitheapResult_bh7_22_c15;
            end if;
            if ce_17 = '1' then
               tmp_bitheapResult_bh7_22_c17 <= tmp_bitheapResult_bh7_22_c16;
            end if;
            if ce_18 = '1' then
               tmp_bitheapResult_bh7_22_c18 <= tmp_bitheapResult_bh7_22_c17;
            end if;
            if ce_19 = '1' then
               tmp_bitheapResult_bh7_22_c19 <= tmp_bitheapResult_bh7_22_c18;
            end if;
            if ce_20 = '1' then
               tmp_bitheapResult_bh7_22_c20 <= tmp_bitheapResult_bh7_22_c19;
            end if;
            if ce_21 = '1' then
               tmp_bitheapResult_bh7_22_c21 <= tmp_bitheapResult_bh7_22_c20;
            end if;
            if ce_22 = '1' then
               tmp_bitheapResult_bh7_22_c22 <= tmp_bitheapResult_bh7_22_c21;
            end if;
            if ce_23 = '1' then
               tmp_bitheapResult_bh7_22_c23 <= tmp_bitheapResult_bh7_22_c22;
            end if;
            if ce_24 = '1' then
               tmp_bitheapResult_bh7_22_c24 <= tmp_bitheapResult_bh7_22_c23;
            end if;
            if ce_25 = '1' then
               tmp_bitheapResult_bh7_22_c25 <= tmp_bitheapResult_bh7_22_c24;
            end if;
            if ce_26 = '1' then
               tmp_bitheapResult_bh7_22_c26 <= tmp_bitheapResult_bh7_22_c25;
            end if;
            if ce_27 = '1' then
               tmp_bitheapResult_bh7_22_c27 <= tmp_bitheapResult_bh7_22_c26;
            end if;
            if ce_28 = '1' then
               tmp_bitheapResult_bh7_22_c28 <= tmp_bitheapResult_bh7_22_c27;
            end if;
            if ce_29 = '1' then
               tmp_bitheapResult_bh7_22_c29 <= tmp_bitheapResult_bh7_22_c28;
            end if;
            if ce_30 = '1' then
               tmp_bitheapResult_bh7_22_c30 <= tmp_bitheapResult_bh7_22_c29;
            end if;
            if ce_31 = '1' then
               tmp_bitheapResult_bh7_22_c31 <= tmp_bitheapResult_bh7_22_c30;
            end if;
            if ce_32 = '1' then
               tmp_bitheapResult_bh7_22_c32 <= tmp_bitheapResult_bh7_22_c31;
            end if;
            if ce_33 = '1' then
               tmp_bitheapResult_bh7_22_c33 <= tmp_bitheapResult_bh7_22_c32;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq800_uid9
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c2);

   tile_0_filtered_output_c2 <= unsigned(tile_0_output_c2(40 downto 0));
   bh7_w0_0_c2 <= tile_0_filtered_output_c2(0);
   bh7_w1_0_c2 <= tile_0_filtered_output_c2(1);
   bh7_w2_0_c2 <= tile_0_filtered_output_c2(2);
   bh7_w3_0_c2 <= tile_0_filtered_output_c2(3);
   bh7_w4_0_c2 <= tile_0_filtered_output_c2(4);
   bh7_w5_0_c2 <= tile_0_filtered_output_c2(5);
   bh7_w6_0_c2 <= tile_0_filtered_output_c2(6);
   bh7_w7_0_c2 <= tile_0_filtered_output_c2(7);
   bh7_w8_0_c2 <= tile_0_filtered_output_c2(8);
   bh7_w9_0_c2 <= tile_0_filtered_output_c2(9);
   bh7_w10_0_c2 <= tile_0_filtered_output_c2(10);
   bh7_w11_0_c2 <= tile_0_filtered_output_c2(11);
   bh7_w12_0_c2 <= tile_0_filtered_output_c2(12);
   bh7_w13_0_c2 <= tile_0_filtered_output_c2(13);
   bh7_w14_0_c2 <= tile_0_filtered_output_c2(14);
   bh7_w15_0_c2 <= tile_0_filtered_output_c2(15);
   bh7_w16_0_c2 <= tile_0_filtered_output_c2(16);
   bh7_w17_0_c2 <= tile_0_filtered_output_c2(17);
   bh7_w18_0_c2 <= tile_0_filtered_output_c2(18);
   bh7_w19_0_c2 <= tile_0_filtered_output_c2(19);
   bh7_w20_0_c2 <= tile_0_filtered_output_c2(20);
   bh7_w21_0_c2 <= tile_0_filtered_output_c2(21);
   bh7_w22_0_c2 <= tile_0_filtered_output_c2(22);
   bh7_w23_0_c2 <= tile_0_filtered_output_c2(23);
   bh7_w24_0_c2 <= tile_0_filtered_output_c2(24);
   bh7_w25_0_c2 <= tile_0_filtered_output_c2(25);
   bh7_w26_0_c2 <= tile_0_filtered_output_c2(26);
   bh7_w27_0_c2 <= tile_0_filtered_output_c2(27);
   bh7_w28_0_c2 <= tile_0_filtered_output_c2(28);
   bh7_w29_0_c2 <= tile_0_filtered_output_c2(29);
   bh7_w30_0_c2 <= tile_0_filtered_output_c2(30);
   bh7_w31_0_c2 <= tile_0_filtered_output_c2(31);
   bh7_w32_0_c2 <= tile_0_filtered_output_c2(32);
   bh7_w33_0_c2 <= tile_0_filtered_output_c2(33);
   bh7_w34_0_c2 <= tile_0_filtered_output_c2(34);
   bh7_w35_0_c2 <= tile_0_filtered_output_c2(35);
   bh7_w36_0_c2 <= tile_0_filtered_output_c2(36);
   bh7_w37_0_c2 <= tile_0_filtered_output_c2(37);
   bh7_w38_0_c2 <= tile_0_filtered_output_c2(38);
   bh7_w39_0_c2 <= tile_0_filtered_output_c2(39);
   bh7_w40_0_c2 <= tile_0_filtered_output_c2(40);
   tile_1_X_c0 <= X(33 downto 17);
   tile_1_Y_c0 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_Freq800_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c2);

   tile_1_filtered_output_c2 <= unsigned(tile_1_output_c2(40 downto 0));
   bh7_w17_1_c2 <= tile_1_filtered_output_c2(0);
   bh7_w18_1_c2 <= tile_1_filtered_output_c2(1);
   bh7_w19_1_c2 <= tile_1_filtered_output_c2(2);
   bh7_w20_1_c2 <= tile_1_filtered_output_c2(3);
   bh7_w21_1_c2 <= tile_1_filtered_output_c2(4);
   bh7_w22_1_c2 <= tile_1_filtered_output_c2(5);
   bh7_w23_1_c2 <= tile_1_filtered_output_c2(6);
   bh7_w24_1_c2 <= tile_1_filtered_output_c2(7);
   bh7_w25_1_c2 <= tile_1_filtered_output_c2(8);
   bh7_w26_1_c2 <= tile_1_filtered_output_c2(9);
   bh7_w27_1_c2 <= tile_1_filtered_output_c2(10);
   bh7_w28_1_c2 <= tile_1_filtered_output_c2(11);
   bh7_w29_1_c2 <= tile_1_filtered_output_c2(12);
   bh7_w30_1_c2 <= tile_1_filtered_output_c2(13);
   bh7_w31_1_c2 <= tile_1_filtered_output_c2(14);
   bh7_w32_1_c2 <= tile_1_filtered_output_c2(15);
   bh7_w33_1_c2 <= tile_1_filtered_output_c2(16);
   bh7_w34_1_c2 <= tile_1_filtered_output_c2(17);
   bh7_w35_1_c2 <= tile_1_filtered_output_c2(18);
   bh7_w36_1_c2 <= tile_1_filtered_output_c2(19);
   bh7_w37_1_c2 <= tile_1_filtered_output_c2(20);
   bh7_w38_1_c2 <= tile_1_filtered_output_c2(21);
   bh7_w39_1_c2 <= tile_1_filtered_output_c2(22);
   bh7_w40_1_c2 <= tile_1_filtered_output_c2(23);
   bh7_w41_0_c2 <= tile_1_filtered_output_c2(24);
   bh7_w42_0_c2 <= tile_1_filtered_output_c2(25);
   bh7_w43_0_c2 <= tile_1_filtered_output_c2(26);
   bh7_w44_0_c2 <= tile_1_filtered_output_c2(27);
   bh7_w45_0_c2 <= tile_1_filtered_output_c2(28);
   bh7_w46_0_c2 <= tile_1_filtered_output_c2(29);
   bh7_w47_0_c2 <= tile_1_filtered_output_c2(30);
   bh7_w48_0_c2 <= tile_1_filtered_output_c2(31);
   bh7_w49_0_c2 <= tile_1_filtered_output_c2(32);
   bh7_w50_0_c2 <= tile_1_filtered_output_c2(33);
   bh7_w51_0_c2 <= tile_1_filtered_output_c2(34);
   bh7_w52_0_c2 <= tile_1_filtered_output_c2(35);
   bh7_w53_0_c2 <= tile_1_filtered_output_c2(36);
   bh7_w54_0_c2 <= tile_1_filtered_output_c2(37);
   bh7_w55_0_c2 <= tile_1_filtered_output_c2(38);
   bh7_w56_0_c2 <= tile_1_filtered_output_c2(39);
   bh7_w57_0_c2 <= tile_1_filtered_output_c2(40);
   tile_2_X_c0 <= X(50 downto 34);
   tile_2_Y_c0 <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_Freq800_uid13
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c2);

   tile_2_filtered_output_c2 <= unsigned(tile_2_output_c2(40 downto 0));
   bh7_w34_2_c2 <= tile_2_filtered_output_c2(0);
   bh7_w35_2_c2 <= tile_2_filtered_output_c2(1);
   bh7_w36_2_c2 <= tile_2_filtered_output_c2(2);
   bh7_w37_2_c2 <= tile_2_filtered_output_c2(3);
   bh7_w38_2_c2 <= tile_2_filtered_output_c2(4);
   bh7_w39_2_c2 <= tile_2_filtered_output_c2(5);
   bh7_w40_2_c2 <= tile_2_filtered_output_c2(6);
   bh7_w41_1_c2 <= tile_2_filtered_output_c2(7);
   bh7_w42_1_c2 <= tile_2_filtered_output_c2(8);
   bh7_w43_1_c2 <= tile_2_filtered_output_c2(9);
   bh7_w44_1_c2 <= tile_2_filtered_output_c2(10);
   bh7_w45_1_c2 <= tile_2_filtered_output_c2(11);
   bh7_w46_1_c2 <= tile_2_filtered_output_c2(12);
   bh7_w47_1_c2 <= tile_2_filtered_output_c2(13);
   bh7_w48_1_c2 <= tile_2_filtered_output_c2(14);
   bh7_w49_1_c2 <= tile_2_filtered_output_c2(15);
   bh7_w50_1_c2 <= tile_2_filtered_output_c2(16);
   bh7_w51_1_c2 <= tile_2_filtered_output_c2(17);
   bh7_w52_1_c2 <= tile_2_filtered_output_c2(18);
   bh7_w53_1_c2 <= tile_2_filtered_output_c2(19);
   bh7_w54_1_c2 <= tile_2_filtered_output_c2(20);
   bh7_w55_1_c2 <= tile_2_filtered_output_c2(21);
   bh7_w56_1_c2 <= tile_2_filtered_output_c2(22);
   bh7_w57_1_c2 <= tile_2_filtered_output_c2(23);
   bh7_w58_0_c2 <= tile_2_filtered_output_c2(24);
   bh7_w59_0_c2 <= tile_2_filtered_output_c2(25);
   bh7_w60_0_c2 <= tile_2_filtered_output_c2(26);
   bh7_w61_0_c2 <= tile_2_filtered_output_c2(27);
   bh7_w62_0_c2 <= tile_2_filtered_output_c2(28);
   bh7_w63_0_c2 <= tile_2_filtered_output_c2(29);
   bh7_w64_0_c2 <= tile_2_filtered_output_c2(30);
   bh7_w65_0_c2 <= tile_2_filtered_output_c2(31);
   bh7_w66_0_c2 <= tile_2_filtered_output_c2(32);
   bh7_w67_0_c2 <= tile_2_filtered_output_c2(33);
   bh7_w68_0_c2 <= tile_2_filtered_output_c2(34);
   bh7_w69_0_c2 <= tile_2_filtered_output_c2(35);
   bh7_w70_0_c2 <= tile_2_filtered_output_c2(36);
   bh7_w71_0_c2 <= tile_2_filtered_output_c2(37);
   bh7_w72_0_c2 <= tile_2_filtered_output_c2(38);
   bh7_w73_0_c2 <= tile_2_filtered_output_c2(39);
   bh7_w74_0_c2 <= tile_2_filtered_output_c2(40);
   tile_3_X_c0 <= X(52 downto 51);
   tile_3_Y_c0 <= Y(23 downto 21);
   tile_3_mult: IntMultiplierLUT_2x3_Freq800_uid15
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w72_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w73_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w74_1_c0 <= tile_3_filtered_output_c0(2);
   bh7_w75_0_c0 <= tile_3_filtered_output_c0(3);
   bh7_w76_0_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(52 downto 51);
   tile_4_Y_c0 <= Y(20 downto 18);
   tile_4_mult: IntMultiplierLUT_2x3_Freq800_uid20
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(4 downto 0));
   bh7_w69_1_c0 <= tile_4_filtered_output_c0(0);
   bh7_w70_1_c0 <= tile_4_filtered_output_c0(1);
   bh7_w71_1_c0 <= tile_4_filtered_output_c0(2);
   bh7_w72_2_c0 <= tile_4_filtered_output_c0(3);
   bh7_w73_2_c0 <= tile_4_filtered_output_c0(4);
   tile_5_X_c0 <= X(52 downto 51);
   tile_5_Y_c0 <= Y(17 downto 15);
   tile_5_mult: IntMultiplierLUT_2x3_Freq800_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w66_1_c0 <= tile_5_filtered_output_c0(0);
   bh7_w67_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w68_1_c0 <= tile_5_filtered_output_c0(2);
   bh7_w69_2_c0 <= tile_5_filtered_output_c0(3);
   bh7_w70_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(52 downto 51);
   tile_6_Y_c0 <= Y(14 downto 12);
   tile_6_mult: IntMultiplierLUT_2x3_Freq800_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w63_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w64_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w65_1_c0 <= tile_6_filtered_output_c0(2);
   bh7_w66_2_c0 <= tile_6_filtered_output_c0(3);
   bh7_w67_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(52 downto 51);
   tile_7_Y_c0 <= Y(11 downto 9);
   tile_7_mult: IntMultiplierLUT_2x3_Freq800_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(4 downto 0));
   bh7_w60_1_c0 <= tile_7_filtered_output_c0(0);
   bh7_w61_1_c0 <= tile_7_filtered_output_c0(1);
   bh7_w62_1_c0 <= tile_7_filtered_output_c0(2);
   bh7_w63_2_c0 <= tile_7_filtered_output_c0(3);
   bh7_w64_2_c0 <= tile_7_filtered_output_c0(4);
   tile_8_X_c0 <= X(52 downto 51);
   tile_8_Y_c0 <= Y(8 downto 6);
   tile_8_mult: IntMultiplierLUT_2x3_Freq800_uid40
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w57_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w58_1_c0 <= tile_8_filtered_output_c0(1);
   bh7_w59_1_c0 <= tile_8_filtered_output_c0(2);
   bh7_w60_2_c0 <= tile_8_filtered_output_c0(3);
   bh7_w61_2_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(52 downto 51);
   tile_9_Y_c0 <= Y(5 downto 3);
   tile_9_mult: IntMultiplierLUT_2x3_Freq800_uid45
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w54_2_c0 <= tile_9_filtered_output_c0(0);
   bh7_w55_2_c0 <= tile_9_filtered_output_c0(1);
   bh7_w56_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w57_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w58_2_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(52 downto 51);
   tile_10_Y_c0 <= Y(2 downto 0);
   tile_10_mult: IntMultiplierLUT_2x3_Freq800_uid50
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(4 downto 0));
   bh7_w51_2_c0 <= tile_10_filtered_output_c0(0);
   bh7_w52_2_c0 <= tile_10_filtered_output_c0(1);
   bh7_w53_2_c0 <= tile_10_filtered_output_c0(2);
   bh7_w54_3_c0 <= tile_10_filtered_output_c0(3);
   bh7_w55_3_c0 <= tile_10_filtered_output_c0(4);
   tile_11_X_c0 <= X(16 downto 0);
   tile_11_Y_c0 <= Y(47 downto 24);
   tile_11_mult: DSPBlock_17x24_Freq800_uid55
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c2);

   tile_11_filtered_output_c2 <= unsigned(tile_11_output_c2(40 downto 0));
   bh7_w24_2_c2 <= tile_11_filtered_output_c2(0);
   bh7_w25_2_c2 <= tile_11_filtered_output_c2(1);
   bh7_w26_2_c2 <= tile_11_filtered_output_c2(2);
   bh7_w27_2_c2 <= tile_11_filtered_output_c2(3);
   bh7_w28_2_c2 <= tile_11_filtered_output_c2(4);
   bh7_w29_2_c2 <= tile_11_filtered_output_c2(5);
   bh7_w30_2_c2 <= tile_11_filtered_output_c2(6);
   bh7_w31_2_c2 <= tile_11_filtered_output_c2(7);
   bh7_w32_2_c2 <= tile_11_filtered_output_c2(8);
   bh7_w33_2_c2 <= tile_11_filtered_output_c2(9);
   bh7_w34_3_c2 <= tile_11_filtered_output_c2(10);
   bh7_w35_3_c2 <= tile_11_filtered_output_c2(11);
   bh7_w36_3_c2 <= tile_11_filtered_output_c2(12);
   bh7_w37_3_c2 <= tile_11_filtered_output_c2(13);
   bh7_w38_3_c2 <= tile_11_filtered_output_c2(14);
   bh7_w39_3_c2 <= tile_11_filtered_output_c2(15);
   bh7_w40_3_c2 <= tile_11_filtered_output_c2(16);
   bh7_w41_2_c2 <= tile_11_filtered_output_c2(17);
   bh7_w42_2_c2 <= tile_11_filtered_output_c2(18);
   bh7_w43_2_c2 <= tile_11_filtered_output_c2(19);
   bh7_w44_2_c2 <= tile_11_filtered_output_c2(20);
   bh7_w45_2_c2 <= tile_11_filtered_output_c2(21);
   bh7_w46_2_c2 <= tile_11_filtered_output_c2(22);
   bh7_w47_2_c2 <= tile_11_filtered_output_c2(23);
   bh7_w48_2_c2 <= tile_11_filtered_output_c2(24);
   bh7_w49_2_c2 <= tile_11_filtered_output_c2(25);
   bh7_w50_2_c2 <= tile_11_filtered_output_c2(26);
   bh7_w51_3_c2 <= tile_11_filtered_output_c2(27);
   bh7_w52_3_c2 <= tile_11_filtered_output_c2(28);
   bh7_w53_3_c2 <= tile_11_filtered_output_c2(29);
   bh7_w54_4_c2 <= tile_11_filtered_output_c2(30);
   bh7_w55_4_c2 <= tile_11_filtered_output_c2(31);
   bh7_w56_3_c2 <= tile_11_filtered_output_c2(32);
   bh7_w57_4_c2 <= tile_11_filtered_output_c2(33);
   bh7_w58_3_c2 <= tile_11_filtered_output_c2(34);
   bh7_w59_2_c2 <= tile_11_filtered_output_c2(35);
   bh7_w60_3_c2 <= tile_11_filtered_output_c2(36);
   bh7_w61_3_c2 <= tile_11_filtered_output_c2(37);
   bh7_w62_2_c2 <= tile_11_filtered_output_c2(38);
   bh7_w63_3_c2 <= tile_11_filtered_output_c2(39);
   bh7_w64_3_c2 <= tile_11_filtered_output_c2(40);
   tile_12_X_c0 <= X(33 downto 17);
   tile_12_Y_c0 <= Y(47 downto 24);
   tile_12_mult: DSPBlock_17x24_Freq800_uid57
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c2);

   tile_12_filtered_output_c2 <= unsigned(tile_12_output_c2(40 downto 0));
   bh7_w41_3_c2 <= tile_12_filtered_output_c2(0);
   bh7_w42_3_c2 <= tile_12_filtered_output_c2(1);
   bh7_w43_3_c2 <= tile_12_filtered_output_c2(2);
   bh7_w44_3_c2 <= tile_12_filtered_output_c2(3);
   bh7_w45_3_c2 <= tile_12_filtered_output_c2(4);
   bh7_w46_3_c2 <= tile_12_filtered_output_c2(5);
   bh7_w47_3_c2 <= tile_12_filtered_output_c2(6);
   bh7_w48_3_c2 <= tile_12_filtered_output_c2(7);
   bh7_w49_3_c2 <= tile_12_filtered_output_c2(8);
   bh7_w50_3_c2 <= tile_12_filtered_output_c2(9);
   bh7_w51_4_c2 <= tile_12_filtered_output_c2(10);
   bh7_w52_4_c2 <= tile_12_filtered_output_c2(11);
   bh7_w53_4_c2 <= tile_12_filtered_output_c2(12);
   bh7_w54_5_c2 <= tile_12_filtered_output_c2(13);
   bh7_w55_5_c2 <= tile_12_filtered_output_c2(14);
   bh7_w56_4_c2 <= tile_12_filtered_output_c2(15);
   bh7_w57_5_c2 <= tile_12_filtered_output_c2(16);
   bh7_w58_4_c2 <= tile_12_filtered_output_c2(17);
   bh7_w59_3_c2 <= tile_12_filtered_output_c2(18);
   bh7_w60_4_c2 <= tile_12_filtered_output_c2(19);
   bh7_w61_4_c2 <= tile_12_filtered_output_c2(20);
   bh7_w62_3_c2 <= tile_12_filtered_output_c2(21);
   bh7_w63_4_c2 <= tile_12_filtered_output_c2(22);
   bh7_w64_4_c2 <= tile_12_filtered_output_c2(23);
   bh7_w65_2_c2 <= tile_12_filtered_output_c2(24);
   bh7_w66_3_c2 <= tile_12_filtered_output_c2(25);
   bh7_w67_3_c2 <= tile_12_filtered_output_c2(26);
   bh7_w68_2_c2 <= tile_12_filtered_output_c2(27);
   bh7_w69_3_c2 <= tile_12_filtered_output_c2(28);
   bh7_w70_3_c2 <= tile_12_filtered_output_c2(29);
   bh7_w71_2_c2 <= tile_12_filtered_output_c2(30);
   bh7_w72_3_c2 <= tile_12_filtered_output_c2(31);
   bh7_w73_3_c2 <= tile_12_filtered_output_c2(32);
   bh7_w74_2_c2 <= tile_12_filtered_output_c2(33);
   bh7_w75_1_c2 <= tile_12_filtered_output_c2(34);
   bh7_w76_1_c2 <= tile_12_filtered_output_c2(35);
   bh7_w77_0_c2 <= tile_12_filtered_output_c2(36);
   bh7_w78_0_c2 <= tile_12_filtered_output_c2(37);
   bh7_w79_0_c2 <= tile_12_filtered_output_c2(38);
   bh7_w80_0_c2 <= tile_12_filtered_output_c2(39);
   bh7_w81_0_c2 <= tile_12_filtered_output_c2(40);
   tile_13_X_c0 <= X(50 downto 34);
   tile_13_Y_c0 <= Y(47 downto 24);
   tile_13_mult: DSPBlock_17x24_Freq800_uid59
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c2);

   tile_13_filtered_output_c2 <= unsigned(tile_13_output_c2(40 downto 0));
   bh7_w58_5_c2 <= tile_13_filtered_output_c2(0);
   bh7_w59_4_c2 <= tile_13_filtered_output_c2(1);
   bh7_w60_5_c2 <= tile_13_filtered_output_c2(2);
   bh7_w61_5_c2 <= tile_13_filtered_output_c2(3);
   bh7_w62_4_c2 <= tile_13_filtered_output_c2(4);
   bh7_w63_5_c2 <= tile_13_filtered_output_c2(5);
   bh7_w64_5_c2 <= tile_13_filtered_output_c2(6);
   bh7_w65_3_c2 <= tile_13_filtered_output_c2(7);
   bh7_w66_4_c2 <= tile_13_filtered_output_c2(8);
   bh7_w67_4_c2 <= tile_13_filtered_output_c2(9);
   bh7_w68_3_c2 <= tile_13_filtered_output_c2(10);
   bh7_w69_4_c2 <= tile_13_filtered_output_c2(11);
   bh7_w70_4_c2 <= tile_13_filtered_output_c2(12);
   bh7_w71_3_c2 <= tile_13_filtered_output_c2(13);
   bh7_w72_4_c2 <= tile_13_filtered_output_c2(14);
   bh7_w73_4_c2 <= tile_13_filtered_output_c2(15);
   bh7_w74_3_c2 <= tile_13_filtered_output_c2(16);
   bh7_w75_2_c2 <= tile_13_filtered_output_c2(17);
   bh7_w76_2_c2 <= tile_13_filtered_output_c2(18);
   bh7_w77_1_c2 <= tile_13_filtered_output_c2(19);
   bh7_w78_1_c2 <= tile_13_filtered_output_c2(20);
   bh7_w79_1_c2 <= tile_13_filtered_output_c2(21);
   bh7_w80_1_c2 <= tile_13_filtered_output_c2(22);
   bh7_w81_1_c2 <= tile_13_filtered_output_c2(23);
   bh7_w82_0_c2 <= tile_13_filtered_output_c2(24);
   bh7_w83_0_c2 <= tile_13_filtered_output_c2(25);
   bh7_w84_0_c2 <= tile_13_filtered_output_c2(26);
   bh7_w85_0_c2 <= tile_13_filtered_output_c2(27);
   bh7_w86_0_c2 <= tile_13_filtered_output_c2(28);
   bh7_w87_0_c2 <= tile_13_filtered_output_c2(29);
   bh7_w88_0_c2 <= tile_13_filtered_output_c2(30);
   bh7_w89_0_c2 <= tile_13_filtered_output_c2(31);
   bh7_w90_0_c2 <= tile_13_filtered_output_c2(32);
   bh7_w91_0_c2 <= tile_13_filtered_output_c2(33);
   bh7_w92_0_c2 <= tile_13_filtered_output_c2(34);
   bh7_w93_0_c2 <= tile_13_filtered_output_c2(35);
   bh7_w94_0_c2 <= tile_13_filtered_output_c2(36);
   bh7_w95_0_c2 <= tile_13_filtered_output_c2(37);
   bh7_w96_0_c2 <= tile_13_filtered_output_c2(38);
   bh7_w97_0_c2 <= tile_13_filtered_output_c2(39);
   bh7_w98_0_c2 <= tile_13_filtered_output_c2(40);
   tile_14_X_c0 <= X(52 downto 51);
   tile_14_Y_c0 <= Y(47 downto 45);
   tile_14_mult: IntMultiplierLUT_2x3_Freq800_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w96_1_c0 <= tile_14_filtered_output_c0(0);
   bh7_w97_1_c0 <= tile_14_filtered_output_c0(1);
   bh7_w98_1_c0 <= tile_14_filtered_output_c0(2);
   bh7_w99_0_c0 <= tile_14_filtered_output_c0(3);
   bh7_w100_0_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(52 downto 51);
   tile_15_Y_c0 <= Y(44 downto 42);
   tile_15_mult: IntMultiplierLUT_2x3_Freq800_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w93_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w94_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w95_1_c0 <= tile_15_filtered_output_c0(2);
   bh7_w96_2_c0 <= tile_15_filtered_output_c0(3);
   bh7_w97_2_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(52 downto 51);
   tile_16_Y_c0 <= Y(41 downto 39);
   tile_16_mult: IntMultiplierLUT_2x3_Freq800_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(4 downto 0));
   bh7_w90_1_c0 <= tile_16_filtered_output_c0(0);
   bh7_w91_1_c0 <= tile_16_filtered_output_c0(1);
   bh7_w92_1_c0 <= tile_16_filtered_output_c0(2);
   bh7_w93_2_c0 <= tile_16_filtered_output_c0(3);
   bh7_w94_2_c0 <= tile_16_filtered_output_c0(4);
   tile_17_X_c0 <= X(52 downto 51);
   tile_17_Y_c0 <= Y(38 downto 36);
   tile_17_mult: IntMultiplierLUT_2x3_Freq800_uid76
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w87_1_c0 <= tile_17_filtered_output_c0(0);
   bh7_w88_1_c0 <= tile_17_filtered_output_c0(1);
   bh7_w89_1_c0 <= tile_17_filtered_output_c0(2);
   bh7_w90_2_c0 <= tile_17_filtered_output_c0(3);
   bh7_w91_2_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(52 downto 51);
   tile_18_Y_c0 <= Y(35 downto 33);
   tile_18_mult: IntMultiplierLUT_2x3_Freq800_uid81
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w84_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w85_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w86_1_c0 <= tile_18_filtered_output_c0(2);
   bh7_w87_2_c0 <= tile_18_filtered_output_c0(3);
   bh7_w88_2_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(52 downto 51);
   tile_19_Y_c0 <= Y(32 downto 30);
   tile_19_mult: IntMultiplierLUT_2x3_Freq800_uid86
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(4 downto 0));
   bh7_w81_2_c0 <= tile_19_filtered_output_c0(0);
   bh7_w82_1_c0 <= tile_19_filtered_output_c0(1);
   bh7_w83_1_c0 <= tile_19_filtered_output_c0(2);
   bh7_w84_2_c0 <= tile_19_filtered_output_c0(3);
   bh7_w85_2_c0 <= tile_19_filtered_output_c0(4);
   tile_20_X_c0 <= X(52 downto 51);
   tile_20_Y_c0 <= Y(29 downto 27);
   tile_20_mult: IntMultiplierLUT_2x3_Freq800_uid91
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w78_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w79_2_c0 <= tile_20_filtered_output_c0(1);
   bh7_w80_2_c0 <= tile_20_filtered_output_c0(2);
   bh7_w81_3_c0 <= tile_20_filtered_output_c0(3);
   bh7_w82_2_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(52 downto 51);
   tile_21_Y_c0 <= Y(26 downto 24);
   tile_21_mult: IntMultiplierLUT_2x3_Freq800_uid96
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w75_3_c0 <= tile_21_filtered_output_c0(0);
   bh7_w76_3_c0 <= tile_21_filtered_output_c0(1);
   bh7_w77_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w78_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w79_3_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(16 downto 16);
   tile_22_Y_c0 <= Y(52 downto 52);
   tile_22_mult: IntMultiplierLUT_1x1_Freq800_uid101
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(0 downto 0));
   bh7_w68_4_c0 <= tile_22_filtered_output_c0(0);
   tile_23_X_c0 <= X(15 downto 12);
   tile_23_Y_c0 <= Y(52 downto 52);
   tile_23_mult: IntMultiplierLUT_4x1_Freq800_uid103
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(3 downto 0));
   bh7_w64_6_c0 <= tile_23_filtered_output_c0(0);
   bh7_w65_4_c0 <= tile_23_filtered_output_c0(1);
   bh7_w66_5_c0 <= tile_23_filtered_output_c0(2);
   bh7_w67_5_c0 <= tile_23_filtered_output_c0(3);
   tile_24_X_c0 <= X(11 downto 8);
   tile_24_Y_c0 <= Y(52 downto 52);
   tile_24_mult: IntMultiplierLUT_4x1_Freq800_uid105
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(3 downto 0));
   bh7_w60_6_c0 <= tile_24_filtered_output_c0(0);
   bh7_w61_6_c0 <= tile_24_filtered_output_c0(1);
   bh7_w62_5_c0 <= tile_24_filtered_output_c0(2);
   bh7_w63_6_c0 <= tile_24_filtered_output_c0(3);
   tile_25_X_c0 <= X(7 downto 4);
   tile_25_Y_c0 <= Y(52 downto 52);
   tile_25_mult: IntMultiplierLUT_4x1_Freq800_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(3 downto 0));
   bh7_w56_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w57_6_c0 <= tile_25_filtered_output_c0(1);
   bh7_w58_6_c0 <= tile_25_filtered_output_c0(2);
   bh7_w59_5_c0 <= tile_25_filtered_output_c0(3);
   tile_26_X_c0 <= X(3 downto 0);
   tile_26_Y_c0 <= Y(52 downto 52);
   tile_26_mult: IntMultiplierLUT_4x1_Freq800_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(3 downto 0));
   bh7_w52_5_c0 <= tile_26_filtered_output_c0(0);
   bh7_w53_5_c0 <= tile_26_filtered_output_c0(1);
   bh7_w54_6_c0 <= tile_26_filtered_output_c0(2);
   bh7_w55_6_c0 <= tile_26_filtered_output_c0(3);
   tile_27_X_c0 <= X(16 downto 15);
   tile_27_Y_c0 <= Y(51 downto 50);
   tile_27_mult: IntMultiplierLUT_2x2_Freq800_uid111
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(3 downto 0));
   bh7_w65_5_c0 <= tile_27_filtered_output_c0(0);
   bh7_w66_6_c0 <= tile_27_filtered_output_c0(1);
   bh7_w67_6_c0 <= tile_27_filtered_output_c0(2);
   bh7_w68_5_c0 <= tile_27_filtered_output_c0(3);
   tile_28_X_c0 <= X(14 downto 12);
   tile_28_Y_c0 <= Y(51 downto 50);
   tile_28_mult: IntMultiplierLUT_3x2_Freq800_uid116
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(4 downto 0));
   bh7_w62_6_c0 <= tile_28_filtered_output_c0(0);
   bh7_w63_7_c0 <= tile_28_filtered_output_c0(1);
   bh7_w64_7_c0 <= tile_28_filtered_output_c0(2);
   bh7_w65_6_c0 <= tile_28_filtered_output_c0(3);
   bh7_w66_7_c0 <= tile_28_filtered_output_c0(4);
   tile_29_X_c0 <= X(11 downto 9);
   tile_29_Y_c0 <= Y(51 downto 50);
   tile_29_mult: IntMultiplierLUT_3x2_Freq800_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w59_6_c0 <= tile_29_filtered_output_c0(0);
   bh7_w60_7_c0 <= tile_29_filtered_output_c0(1);
   bh7_w61_7_c0 <= tile_29_filtered_output_c0(2);
   bh7_w62_7_c0 <= tile_29_filtered_output_c0(3);
   bh7_w63_8_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(8 downto 6);
   tile_30_Y_c0 <= Y(51 downto 50);
   tile_30_mult: IntMultiplierLUT_3x2_Freq800_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w56_6_c0 <= tile_30_filtered_output_c0(0);
   bh7_w57_7_c0 <= tile_30_filtered_output_c0(1);
   bh7_w58_7_c0 <= tile_30_filtered_output_c0(2);
   bh7_w59_7_c0 <= tile_30_filtered_output_c0(3);
   bh7_w60_8_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(5 downto 3);
   tile_31_Y_c0 <= Y(51 downto 50);
   tile_31_mult: IntMultiplierLUT_3x2_Freq800_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(4 downto 0));
   bh7_w53_6_c0 <= tile_31_filtered_output_c0(0);
   bh7_w54_7_c0 <= tile_31_filtered_output_c0(1);
   bh7_w55_7_c0 <= tile_31_filtered_output_c0(2);
   bh7_w56_7_c0 <= tile_31_filtered_output_c0(3);
   bh7_w57_8_c0 <= tile_31_filtered_output_c0(4);
   tile_32_X_c0 <= X(2 downto 0);
   tile_32_Y_c0 <= Y(51 downto 50);
   tile_32_mult: IntMultiplierLUT_3x2_Freq800_uid136
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w50_4_c0 <= tile_32_filtered_output_c0(0);
   bh7_w51_5_c0 <= tile_32_filtered_output_c0(1);
   bh7_w52_6_c0 <= tile_32_filtered_output_c0(2);
   bh7_w53_7_c0 <= tile_32_filtered_output_c0(3);
   bh7_w54_8_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(16 downto 15);
   tile_33_Y_c0 <= Y(49 downto 48);
   tile_33_mult: IntMultiplierLUT_2x2_Freq800_uid141
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(3 downto 0));
   bh7_w63_9_c0 <= tile_33_filtered_output_c0(0);
   bh7_w64_8_c0 <= tile_33_filtered_output_c0(1);
   bh7_w65_7_c0 <= tile_33_filtered_output_c0(2);
   bh7_w66_8_c0 <= tile_33_filtered_output_c0(3);
   tile_34_X_c0 <= X(14 downto 12);
   tile_34_Y_c0 <= Y(49 downto 48);
   tile_34_mult: IntMultiplierLUT_3x2_Freq800_uid146
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(4 downto 0));
   bh7_w60_9_c0 <= tile_34_filtered_output_c0(0);
   bh7_w61_8_c0 <= tile_34_filtered_output_c0(1);
   bh7_w62_8_c0 <= tile_34_filtered_output_c0(2);
   bh7_w63_10_c0 <= tile_34_filtered_output_c0(3);
   bh7_w64_9_c0 <= tile_34_filtered_output_c0(4);
   tile_35_X_c0 <= X(11 downto 9);
   tile_35_Y_c0 <= Y(49 downto 48);
   tile_35_mult: IntMultiplierLUT_3x2_Freq800_uid151
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w57_9_c0 <= tile_35_filtered_output_c0(0);
   bh7_w58_8_c0 <= tile_35_filtered_output_c0(1);
   bh7_w59_8_c0 <= tile_35_filtered_output_c0(2);
   bh7_w60_10_c0 <= tile_35_filtered_output_c0(3);
   bh7_w61_9_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(8 downto 6);
   tile_36_Y_c0 <= Y(49 downto 48);
   tile_36_mult: IntMultiplierLUT_3x2_Freq800_uid156
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w54_9_c0 <= tile_36_filtered_output_c0(0);
   bh7_w55_8_c0 <= tile_36_filtered_output_c0(1);
   bh7_w56_8_c0 <= tile_36_filtered_output_c0(2);
   bh7_w57_10_c0 <= tile_36_filtered_output_c0(3);
   bh7_w58_9_c0 <= tile_36_filtered_output_c0(4);
   tile_37_X_c0 <= X(5 downto 3);
   tile_37_Y_c0 <= Y(49 downto 48);
   tile_37_mult: IntMultiplierLUT_3x2_Freq800_uid161
      port map ( clk  => clk,
                 X => tile_37_X_c0,
                 Y => tile_37_Y_c0,
                 R => tile_37_output_c0);

   tile_37_filtered_output_c0 <= unsigned(tile_37_output_c0(4 downto 0));
   bh7_w51_6_c0 <= tile_37_filtered_output_c0(0);
   bh7_w52_7_c0 <= tile_37_filtered_output_c0(1);
   bh7_w53_8_c0 <= tile_37_filtered_output_c0(2);
   bh7_w54_10_c0 <= tile_37_filtered_output_c0(3);
   bh7_w55_9_c0 <= tile_37_filtered_output_c0(4);
   tile_38_X_c0 <= X(2 downto 0);
   tile_38_Y_c0 <= Y(49 downto 48);
   tile_38_mult: IntMultiplierLUT_3x2_Freq800_uid166
      port map ( clk  => clk,
                 X => tile_38_X_c0,
                 Y => tile_38_Y_c0,
                 R => tile_38_output_c0);

   tile_38_filtered_output_c0 <= unsigned(tile_38_output_c0(4 downto 0));
   bh7_w48_4_c0 <= tile_38_filtered_output_c0(0);
   bh7_w49_4_c0 <= tile_38_filtered_output_c0(1);
   bh7_w50_5_c0 <= tile_38_filtered_output_c0(2);
   bh7_w51_7_c0 <= tile_38_filtered_output_c0(3);
   bh7_w52_8_c0 <= tile_38_filtered_output_c0(4);
   tile_39_X_c0 <= X(33 downto 33);
   tile_39_Y_c0 <= Y(52 downto 52);
   tile_39_mult: IntMultiplierLUT_1x1_Freq800_uid171
      port map ( clk  => clk,
                 X => tile_39_X_c0,
                 Y => tile_39_Y_c0,
                 R => tile_39_output_c0);

   tile_39_filtered_output_c0 <= unsigned(tile_39_output_c0(0 downto 0));
   bh7_w85_3_c0 <= tile_39_filtered_output_c0(0);
   tile_40_X_c0 <= X(32 downto 29);
   tile_40_Y_c0 <= Y(52 downto 52);
   tile_40_mult: IntMultiplierLUT_4x1_Freq800_uid173
      port map ( clk  => clk,
                 X => tile_40_X_c0,
                 Y => tile_40_Y_c0,
                 R => tile_40_output_c0);

   tile_40_filtered_output_c0 <= unsigned(tile_40_output_c0(3 downto 0));
   bh7_w81_4_c0 <= tile_40_filtered_output_c0(0);
   bh7_w82_3_c0 <= tile_40_filtered_output_c0(1);
   bh7_w83_2_c0 <= tile_40_filtered_output_c0(2);
   bh7_w84_3_c0 <= tile_40_filtered_output_c0(3);
   tile_41_X_c0 <= X(28 downto 25);
   tile_41_Y_c0 <= Y(52 downto 52);
   tile_41_mult: IntMultiplierLUT_4x1_Freq800_uid175
      port map ( clk  => clk,
                 X => tile_41_X_c0,
                 Y => tile_41_Y_c0,
                 R => tile_41_output_c0);

   tile_41_filtered_output_c0 <= unsigned(tile_41_output_c0(3 downto 0));
   bh7_w77_3_c0 <= tile_41_filtered_output_c0(0);
   bh7_w78_4_c0 <= tile_41_filtered_output_c0(1);
   bh7_w79_4_c0 <= tile_41_filtered_output_c0(2);
   bh7_w80_3_c0 <= tile_41_filtered_output_c0(3);
   tile_42_X_c0 <= X(24 downto 21);
   tile_42_Y_c0 <= Y(52 downto 52);
   tile_42_mult: IntMultiplierLUT_4x1_Freq800_uid177
      port map ( clk  => clk,
                 X => tile_42_X_c0,
                 Y => tile_42_Y_c0,
                 R => tile_42_output_c0);

   tile_42_filtered_output_c0 <= unsigned(tile_42_output_c0(3 downto 0));
   bh7_w73_5_c0 <= tile_42_filtered_output_c0(0);
   bh7_w74_4_c0 <= tile_42_filtered_output_c0(1);
   bh7_w75_4_c0 <= tile_42_filtered_output_c0(2);
   bh7_w76_4_c0 <= tile_42_filtered_output_c0(3);
   tile_43_X_c0 <= X(20 downto 17);
   tile_43_Y_c0 <= Y(52 downto 52);
   tile_43_mult: IntMultiplierLUT_4x1_Freq800_uid179
      port map ( clk  => clk,
                 X => tile_43_X_c0,
                 Y => tile_43_Y_c0,
                 R => tile_43_output_c0);

   tile_43_filtered_output_c0 <= unsigned(tile_43_output_c0(3 downto 0));
   bh7_w69_5_c0 <= tile_43_filtered_output_c0(0);
   bh7_w70_5_c0 <= tile_43_filtered_output_c0(1);
   bh7_w71_4_c0 <= tile_43_filtered_output_c0(2);
   bh7_w72_5_c0 <= tile_43_filtered_output_c0(3);
   tile_44_X_c0 <= X(33 downto 32);
   tile_44_Y_c0 <= Y(51 downto 50);
   tile_44_mult: IntMultiplierLUT_2x2_Freq800_uid181
      port map ( clk  => clk,
                 X => tile_44_X_c0,
                 Y => tile_44_Y_c0,
                 R => tile_44_output_c0);

   tile_44_filtered_output_c0 <= unsigned(tile_44_output_c0(3 downto 0));
   bh7_w82_4_c0 <= tile_44_filtered_output_c0(0);
   bh7_w83_3_c0 <= tile_44_filtered_output_c0(1);
   bh7_w84_4_c0 <= tile_44_filtered_output_c0(2);
   bh7_w85_4_c0 <= tile_44_filtered_output_c0(3);
   tile_45_X_c0 <= X(31 downto 29);
   tile_45_Y_c0 <= Y(51 downto 50);
   tile_45_mult: IntMultiplierLUT_3x2_Freq800_uid186
      port map ( clk  => clk,
                 X => tile_45_X_c0,
                 Y => tile_45_Y_c0,
                 R => tile_45_output_c0);

   tile_45_filtered_output_c0 <= unsigned(tile_45_output_c0(4 downto 0));
   bh7_w79_5_c0 <= tile_45_filtered_output_c0(0);
   bh7_w80_4_c0 <= tile_45_filtered_output_c0(1);
   bh7_w81_5_c0 <= tile_45_filtered_output_c0(2);
   bh7_w82_5_c0 <= tile_45_filtered_output_c0(3);
   bh7_w83_4_c0 <= tile_45_filtered_output_c0(4);
   tile_46_X_c0 <= X(28 downto 26);
   tile_46_Y_c0 <= Y(51 downto 50);
   tile_46_mult: IntMultiplierLUT_3x2_Freq800_uid191
      port map ( clk  => clk,
                 X => tile_46_X_c0,
                 Y => tile_46_Y_c0,
                 R => tile_46_output_c0);

   tile_46_filtered_output_c0 <= unsigned(tile_46_output_c0(4 downto 0));
   bh7_w76_5_c0 <= tile_46_filtered_output_c0(0);
   bh7_w77_4_c0 <= tile_46_filtered_output_c0(1);
   bh7_w78_5_c0 <= tile_46_filtered_output_c0(2);
   bh7_w79_6_c0 <= tile_46_filtered_output_c0(3);
   bh7_w80_5_c0 <= tile_46_filtered_output_c0(4);
   tile_47_X_c0 <= X(25 downto 23);
   tile_47_Y_c0 <= Y(51 downto 50);
   tile_47_mult: IntMultiplierLUT_3x2_Freq800_uid196
      port map ( clk  => clk,
                 X => tile_47_X_c0,
                 Y => tile_47_Y_c0,
                 R => tile_47_output_c0);

   tile_47_filtered_output_c0 <= unsigned(tile_47_output_c0(4 downto 0));
   bh7_w73_6_c0 <= tile_47_filtered_output_c0(0);
   bh7_w74_5_c0 <= tile_47_filtered_output_c0(1);
   bh7_w75_5_c0 <= tile_47_filtered_output_c0(2);
   bh7_w76_6_c0 <= tile_47_filtered_output_c0(3);
   bh7_w77_5_c0 <= tile_47_filtered_output_c0(4);
   tile_48_X_c0 <= X(22 downto 20);
   tile_48_Y_c0 <= Y(51 downto 50);
   tile_48_mult: IntMultiplierLUT_3x2_Freq800_uid201
      port map ( clk  => clk,
                 X => tile_48_X_c0,
                 Y => tile_48_Y_c0,
                 R => tile_48_output_c0);

   tile_48_filtered_output_c0 <= unsigned(tile_48_output_c0(4 downto 0));
   bh7_w70_6_c0 <= tile_48_filtered_output_c0(0);
   bh7_w71_5_c0 <= tile_48_filtered_output_c0(1);
   bh7_w72_6_c0 <= tile_48_filtered_output_c0(2);
   bh7_w73_7_c0 <= tile_48_filtered_output_c0(3);
   bh7_w74_6_c0 <= tile_48_filtered_output_c0(4);
   tile_49_X_c0 <= X(19 downto 17);
   tile_49_Y_c0 <= Y(51 downto 50);
   tile_49_mult: IntMultiplierLUT_3x2_Freq800_uid206
      port map ( clk  => clk,
                 X => tile_49_X_c0,
                 Y => tile_49_Y_c0,
                 R => tile_49_output_c0);

   tile_49_filtered_output_c0 <= unsigned(tile_49_output_c0(4 downto 0));
   bh7_w67_7_c0 <= tile_49_filtered_output_c0(0);
   bh7_w68_6_c0 <= tile_49_filtered_output_c0(1);
   bh7_w69_6_c0 <= tile_49_filtered_output_c0(2);
   bh7_w70_7_c0 <= tile_49_filtered_output_c0(3);
   bh7_w71_6_c0 <= tile_49_filtered_output_c0(4);
   tile_50_X_c0 <= X(33 downto 32);
   tile_50_Y_c0 <= Y(49 downto 48);
   tile_50_mult: IntMultiplierLUT_2x2_Freq800_uid211
      port map ( clk  => clk,
                 X => tile_50_X_c0,
                 Y => tile_50_Y_c0,
                 R => tile_50_output_c0);

   tile_50_filtered_output_c0 <= unsigned(tile_50_output_c0(3 downto 0));
   bh7_w80_6_c0 <= tile_50_filtered_output_c0(0);
   bh7_w81_6_c0 <= tile_50_filtered_output_c0(1);
   bh7_w82_6_c0 <= tile_50_filtered_output_c0(2);
   bh7_w83_5_c0 <= tile_50_filtered_output_c0(3);
   tile_51_X_c0 <= X(31 downto 29);
   tile_51_Y_c0 <= Y(49 downto 48);
   tile_51_mult: IntMultiplierLUT_3x2_Freq800_uid216
      port map ( clk  => clk,
                 X => tile_51_X_c0,
                 Y => tile_51_Y_c0,
                 R => tile_51_output_c0);

   tile_51_filtered_output_c0 <= unsigned(tile_51_output_c0(4 downto 0));
   bh7_w77_6_c0 <= tile_51_filtered_output_c0(0);
   bh7_w78_6_c0 <= tile_51_filtered_output_c0(1);
   bh7_w79_7_c0 <= tile_51_filtered_output_c0(2);
   bh7_w80_7_c0 <= tile_51_filtered_output_c0(3);
   bh7_w81_7_c0 <= tile_51_filtered_output_c0(4);
   tile_52_X_c0 <= X(28 downto 26);
   tile_52_Y_c0 <= Y(49 downto 48);
   tile_52_mult: IntMultiplierLUT_3x2_Freq800_uid221
      port map ( clk  => clk,
                 X => tile_52_X_c0,
                 Y => tile_52_Y_c0,
                 R => tile_52_output_c0);

   tile_52_filtered_output_c0 <= unsigned(tile_52_output_c0(4 downto 0));
   bh7_w74_7_c0 <= tile_52_filtered_output_c0(0);
   bh7_w75_6_c0 <= tile_52_filtered_output_c0(1);
   bh7_w76_7_c0 <= tile_52_filtered_output_c0(2);
   bh7_w77_7_c0 <= tile_52_filtered_output_c0(3);
   bh7_w78_7_c0 <= tile_52_filtered_output_c0(4);
   tile_53_X_c0 <= X(25 downto 23);
   tile_53_Y_c0 <= Y(49 downto 48);
   tile_53_mult: IntMultiplierLUT_3x2_Freq800_uid226
      port map ( clk  => clk,
                 X => tile_53_X_c0,
                 Y => tile_53_Y_c0,
                 R => tile_53_output_c0);

   tile_53_filtered_output_c0 <= unsigned(tile_53_output_c0(4 downto 0));
   bh7_w71_7_c0 <= tile_53_filtered_output_c0(0);
   bh7_w72_7_c0 <= tile_53_filtered_output_c0(1);
   bh7_w73_8_c0 <= tile_53_filtered_output_c0(2);
   bh7_w74_8_c0 <= tile_53_filtered_output_c0(3);
   bh7_w75_7_c0 <= tile_53_filtered_output_c0(4);
   tile_54_X_c0 <= X(22 downto 20);
   tile_54_Y_c0 <= Y(49 downto 48);
   tile_54_mult: IntMultiplierLUT_3x2_Freq800_uid231
      port map ( clk  => clk,
                 X => tile_54_X_c0,
                 Y => tile_54_Y_c0,
                 R => tile_54_output_c0);

   tile_54_filtered_output_c0 <= unsigned(tile_54_output_c0(4 downto 0));
   bh7_w68_7_c0 <= tile_54_filtered_output_c0(0);
   bh7_w69_7_c0 <= tile_54_filtered_output_c0(1);
   bh7_w70_8_c0 <= tile_54_filtered_output_c0(2);
   bh7_w71_8_c0 <= tile_54_filtered_output_c0(3);
   bh7_w72_8_c0 <= tile_54_filtered_output_c0(4);
   tile_55_X_c0 <= X(19 downto 17);
   tile_55_Y_c0 <= Y(49 downto 48);
   tile_55_mult: IntMultiplierLUT_3x2_Freq800_uid236
      port map ( clk  => clk,
                 X => tile_55_X_c0,
                 Y => tile_55_Y_c0,
                 R => tile_55_output_c0);

   tile_55_filtered_output_c0 <= unsigned(tile_55_output_c0(4 downto 0));
   bh7_w65_8_c0 <= tile_55_filtered_output_c0(0);
   bh7_w66_9_c0 <= tile_55_filtered_output_c0(1);
   bh7_w67_8_c0 <= tile_55_filtered_output_c0(2);
   bh7_w68_8_c0 <= tile_55_filtered_output_c0(3);
   bh7_w69_8_c0 <= tile_55_filtered_output_c0(4);
   tile_56_X_c0 <= X(50 downto 50);
   tile_56_Y_c0 <= Y(52 downto 52);
   tile_56_mult: IntMultiplierLUT_1x1_Freq800_uid241
      port map ( clk  => clk,
                 X => tile_56_X_c0,
                 Y => tile_56_Y_c0,
                 R => tile_56_output_c0);

   tile_56_filtered_output_c0 <= unsigned(tile_56_output_c0(0 downto 0));
   bh7_w102_0_c0 <= tile_56_filtered_output_c0(0);
   tile_57_X_c0 <= X(49 downto 46);
   tile_57_Y_c0 <= Y(52 downto 52);
   tile_57_mult: IntMultiplierLUT_4x1_Freq800_uid243
      port map ( clk  => clk,
                 X => tile_57_X_c0,
                 Y => tile_57_Y_c0,
                 R => tile_57_output_c0);

   tile_57_filtered_output_c0 <= unsigned(tile_57_output_c0(3 downto 0));
   bh7_w98_2_c0 <= tile_57_filtered_output_c0(0);
   bh7_w99_1_c0 <= tile_57_filtered_output_c0(1);
   bh7_w100_1_c0 <= tile_57_filtered_output_c0(2);
   bh7_w101_0_c0 <= tile_57_filtered_output_c0(3);
   tile_58_X_c0 <= X(45 downto 42);
   tile_58_Y_c0 <= Y(52 downto 52);
   tile_58_mult: IntMultiplierLUT_4x1_Freq800_uid245
      port map ( clk  => clk,
                 X => tile_58_X_c0,
                 Y => tile_58_Y_c0,
                 R => tile_58_output_c0);

   tile_58_filtered_output_c0 <= unsigned(tile_58_output_c0(3 downto 0));
   bh7_w94_3_c0 <= tile_58_filtered_output_c0(0);
   bh7_w95_2_c0 <= tile_58_filtered_output_c0(1);
   bh7_w96_3_c0 <= tile_58_filtered_output_c0(2);
   bh7_w97_3_c0 <= tile_58_filtered_output_c0(3);
   tile_59_X_c0 <= X(41 downto 38);
   tile_59_Y_c0 <= Y(52 downto 52);
   tile_59_mult: IntMultiplierLUT_4x1_Freq800_uid247
      port map ( clk  => clk,
                 X => tile_59_X_c0,
                 Y => tile_59_Y_c0,
                 R => tile_59_output_c0);

   tile_59_filtered_output_c0 <= unsigned(tile_59_output_c0(3 downto 0));
   bh7_w90_3_c0 <= tile_59_filtered_output_c0(0);
   bh7_w91_3_c0 <= tile_59_filtered_output_c0(1);
   bh7_w92_2_c0 <= tile_59_filtered_output_c0(2);
   bh7_w93_3_c0 <= tile_59_filtered_output_c0(3);
   tile_60_X_c0 <= X(37 downto 34);
   tile_60_Y_c0 <= Y(52 downto 52);
   tile_60_mult: IntMultiplierLUT_4x1_Freq800_uid249
      port map ( clk  => clk,
                 X => tile_60_X_c0,
                 Y => tile_60_Y_c0,
                 R => tile_60_output_c0);

   tile_60_filtered_output_c0 <= unsigned(tile_60_output_c0(3 downto 0));
   bh7_w86_2_c0 <= tile_60_filtered_output_c0(0);
   bh7_w87_3_c0 <= tile_60_filtered_output_c0(1);
   bh7_w88_3_c0 <= tile_60_filtered_output_c0(2);
   bh7_w89_2_c0 <= tile_60_filtered_output_c0(3);
   tile_61_X_c0 <= X(50 downto 49);
   tile_61_Y_c0 <= Y(51 downto 50);
   tile_61_mult: IntMultiplierLUT_2x2_Freq800_uid251
      port map ( clk  => clk,
                 X => tile_61_X_c0,
                 Y => tile_61_Y_c0,
                 R => tile_61_output_c0);

   tile_61_filtered_output_c0 <= unsigned(tile_61_output_c0(3 downto 0));
   bh7_w99_2_c0 <= tile_61_filtered_output_c0(0);
   bh7_w100_2_c0 <= tile_61_filtered_output_c0(1);
   bh7_w101_1_c0 <= tile_61_filtered_output_c0(2);
   bh7_w102_1_c0 <= tile_61_filtered_output_c0(3);
   tile_62_X_c0 <= X(48 downto 46);
   tile_62_Y_c0 <= Y(51 downto 50);
   tile_62_mult: IntMultiplierLUT_3x2_Freq800_uid256
      port map ( clk  => clk,
                 X => tile_62_X_c0,
                 Y => tile_62_Y_c0,
                 R => tile_62_output_c0);

   tile_62_filtered_output_c0 <= unsigned(tile_62_output_c0(4 downto 0));
   bh7_w96_4_c0 <= tile_62_filtered_output_c0(0);
   bh7_w97_4_c0 <= tile_62_filtered_output_c0(1);
   bh7_w98_3_c0 <= tile_62_filtered_output_c0(2);
   bh7_w99_3_c0 <= tile_62_filtered_output_c0(3);
   bh7_w100_3_c0 <= tile_62_filtered_output_c0(4);
   tile_63_X_c0 <= X(45 downto 43);
   tile_63_Y_c0 <= Y(51 downto 50);
   tile_63_mult: IntMultiplierLUT_3x2_Freq800_uid261
      port map ( clk  => clk,
                 X => tile_63_X_c0,
                 Y => tile_63_Y_c0,
                 R => tile_63_output_c0);

   tile_63_filtered_output_c0 <= unsigned(tile_63_output_c0(4 downto 0));
   bh7_w93_4_c0 <= tile_63_filtered_output_c0(0);
   bh7_w94_4_c0 <= tile_63_filtered_output_c0(1);
   bh7_w95_3_c0 <= tile_63_filtered_output_c0(2);
   bh7_w96_5_c0 <= tile_63_filtered_output_c0(3);
   bh7_w97_5_c0 <= tile_63_filtered_output_c0(4);
   tile_64_X_c0 <= X(42 downto 40);
   tile_64_Y_c0 <= Y(51 downto 50);
   tile_64_mult: IntMultiplierLUT_3x2_Freq800_uid266
      port map ( clk  => clk,
                 X => tile_64_X_c0,
                 Y => tile_64_Y_c0,
                 R => tile_64_output_c0);

   tile_64_filtered_output_c0 <= unsigned(tile_64_output_c0(4 downto 0));
   bh7_w90_4_c0 <= tile_64_filtered_output_c0(0);
   bh7_w91_4_c0 <= tile_64_filtered_output_c0(1);
   bh7_w92_3_c0 <= tile_64_filtered_output_c0(2);
   bh7_w93_5_c0 <= tile_64_filtered_output_c0(3);
   bh7_w94_5_c0 <= tile_64_filtered_output_c0(4);
   tile_65_X_c0 <= X(39 downto 37);
   tile_65_Y_c0 <= Y(51 downto 50);
   tile_65_mult: IntMultiplierLUT_3x2_Freq800_uid271
      port map ( clk  => clk,
                 X => tile_65_X_c0,
                 Y => tile_65_Y_c0,
                 R => tile_65_output_c0);

   tile_65_filtered_output_c0 <= unsigned(tile_65_output_c0(4 downto 0));
   bh7_w87_4_c0 <= tile_65_filtered_output_c0(0);
   bh7_w88_4_c0 <= tile_65_filtered_output_c0(1);
   bh7_w89_3_c0 <= tile_65_filtered_output_c0(2);
   bh7_w90_5_c0 <= tile_65_filtered_output_c0(3);
   bh7_w91_5_c0 <= tile_65_filtered_output_c0(4);
   tile_66_X_c0 <= X(36 downto 34);
   tile_66_Y_c0 <= Y(51 downto 50);
   tile_66_mult: IntMultiplierLUT_3x2_Freq800_uid276
      port map ( clk  => clk,
                 X => tile_66_X_c0,
                 Y => tile_66_Y_c0,
                 R => tile_66_output_c0);

   tile_66_filtered_output_c0 <= unsigned(tile_66_output_c0(4 downto 0));
   bh7_w84_5_c0 <= tile_66_filtered_output_c0(0);
   bh7_w85_5_c0 <= tile_66_filtered_output_c0(1);
   bh7_w86_3_c0 <= tile_66_filtered_output_c0(2);
   bh7_w87_5_c0 <= tile_66_filtered_output_c0(3);
   bh7_w88_5_c0 <= tile_66_filtered_output_c0(4);
   tile_67_X_c0 <= X(50 downto 49);
   tile_67_Y_c0 <= Y(49 downto 48);
   tile_67_mult: IntMultiplierLUT_2x2_Freq800_uid281
      port map ( clk  => clk,
                 X => tile_67_X_c0,
                 Y => tile_67_Y_c0,
                 R => tile_67_output_c0);

   tile_67_filtered_output_c0 <= unsigned(tile_67_output_c0(3 downto 0));
   bh7_w97_6_c0 <= tile_67_filtered_output_c0(0);
   bh7_w98_4_c0 <= tile_67_filtered_output_c0(1);
   bh7_w99_4_c0 <= tile_67_filtered_output_c0(2);
   bh7_w100_4_c0 <= tile_67_filtered_output_c0(3);
   tile_68_X_c0 <= X(48 downto 46);
   tile_68_Y_c0 <= Y(49 downto 48);
   tile_68_mult: IntMultiplierLUT_3x2_Freq800_uid286
      port map ( clk  => clk,
                 X => tile_68_X_c0,
                 Y => tile_68_Y_c0,
                 R => tile_68_output_c0);

   tile_68_filtered_output_c0 <= unsigned(tile_68_output_c0(4 downto 0));
   bh7_w94_6_c0 <= tile_68_filtered_output_c0(0);
   bh7_w95_4_c0 <= tile_68_filtered_output_c0(1);
   bh7_w96_6_c0 <= tile_68_filtered_output_c0(2);
   bh7_w97_7_c0 <= tile_68_filtered_output_c0(3);
   bh7_w98_5_c0 <= tile_68_filtered_output_c0(4);
   tile_69_X_c0 <= X(45 downto 43);
   tile_69_Y_c0 <= Y(49 downto 48);
   tile_69_mult: IntMultiplierLUT_3x2_Freq800_uid291
      port map ( clk  => clk,
                 X => tile_69_X_c0,
                 Y => tile_69_Y_c0,
                 R => tile_69_output_c0);

   tile_69_filtered_output_c0 <= unsigned(tile_69_output_c0(4 downto 0));
   bh7_w91_6_c0 <= tile_69_filtered_output_c0(0);
   bh7_w92_4_c0 <= tile_69_filtered_output_c0(1);
   bh7_w93_6_c0 <= tile_69_filtered_output_c0(2);
   bh7_w94_7_c0 <= tile_69_filtered_output_c0(3);
   bh7_w95_5_c0 <= tile_69_filtered_output_c0(4);
   tile_70_X_c0 <= X(42 downto 40);
   tile_70_Y_c0 <= Y(49 downto 48);
   tile_70_mult: IntMultiplierLUT_3x2_Freq800_uid296
      port map ( clk  => clk,
                 X => tile_70_X_c0,
                 Y => tile_70_Y_c0,
                 R => tile_70_output_c0);

   tile_70_filtered_output_c0 <= unsigned(tile_70_output_c0(4 downto 0));
   bh7_w88_6_c0 <= tile_70_filtered_output_c0(0);
   bh7_w89_4_c0 <= tile_70_filtered_output_c0(1);
   bh7_w90_6_c0 <= tile_70_filtered_output_c0(2);
   bh7_w91_7_c0 <= tile_70_filtered_output_c0(3);
   bh7_w92_5_c0 <= tile_70_filtered_output_c0(4);
   tile_71_X_c0 <= X(39 downto 37);
   tile_71_Y_c0 <= Y(49 downto 48);
   tile_71_mult: IntMultiplierLUT_3x2_Freq800_uid301
      port map ( clk  => clk,
                 X => tile_71_X_c0,
                 Y => tile_71_Y_c0,
                 R => tile_71_output_c0);

   tile_71_filtered_output_c0 <= unsigned(tile_71_output_c0(4 downto 0));
   bh7_w85_6_c0 <= tile_71_filtered_output_c0(0);
   bh7_w86_4_c0 <= tile_71_filtered_output_c0(1);
   bh7_w87_6_c0 <= tile_71_filtered_output_c0(2);
   bh7_w88_7_c0 <= tile_71_filtered_output_c0(3);
   bh7_w89_5_c0 <= tile_71_filtered_output_c0(4);
   tile_72_X_c0 <= X(36 downto 34);
   tile_72_Y_c0 <= Y(49 downto 48);
   tile_72_mult: IntMultiplierLUT_3x2_Freq800_uid306
      port map ( clk  => clk,
                 X => tile_72_X_c0,
                 Y => tile_72_Y_c0,
                 R => tile_72_output_c0);

   tile_72_filtered_output_c0 <= unsigned(tile_72_output_c0(4 downto 0));
   bh7_w82_7_c0 <= tile_72_filtered_output_c0(0);
   bh7_w83_6_c0 <= tile_72_filtered_output_c0(1);
   bh7_w84_6_c0 <= tile_72_filtered_output_c0(2);
   bh7_w85_7_c0 <= tile_72_filtered_output_c0(3);
   bh7_w86_5_c0 <= tile_72_filtered_output_c0(4);
   tile_73_X_c0 <= X(52 downto 51);
   tile_73_Y_c0 <= Y(52 downto 51);
   tile_73_mult: IntMultiplierLUT_2x2_Freq800_uid311
      port map ( clk  => clk,
                 X => tile_73_X_c0,
                 Y => tile_73_Y_c0,
                 R => tile_73_output_c0);

   tile_73_filtered_output_c0 <= unsigned(tile_73_output_c0(3 downto 0));
   bh7_w102_2_c0 <= tile_73_filtered_output_c0(0);
   bh7_w103_0_c0 <= tile_73_filtered_output_c0(1);
   bh7_w104_0_c0 <= tile_73_filtered_output_c0(2);
   bh7_w105_0_c0 <= tile_73_filtered_output_c0(3);
   tile_74_X_c0 <= X(52 downto 51);
   tile_74_Y_c0 <= Y(50 downto 48);
   tile_74_mult: IntMultiplierLUT_2x3_Freq800_uid316
      port map ( clk  => clk,
                 X => tile_74_X_c0,
                 Y => tile_74_Y_c0,
                 R => tile_74_output_c0);

   tile_74_filtered_output_c0 <= unsigned(tile_74_output_c0(4 downto 0));
   bh7_w99_5_c0 <= tile_74_filtered_output_c0(0);
   bh7_w100_5_c0 <= tile_74_filtered_output_c0(1);
   bh7_w101_2_c0 <= tile_74_filtered_output_c0(2);
   bh7_w102_3_c0 <= tile_74_filtered_output_c0(3);
   bh7_w103_1_c0 <= tile_74_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq800_uid322_bh7_uid323_In0_c0 <= "" & bh7_w49_4_c0 & "0" & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid323_In1_c0 <= "" & bh7_w50_4_c0 & bh7_w50_5_c0;
   bh7_w49_5_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1(0);
   bh7_w50_6_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1(1);
   bh7_w51_8_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid323: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid323_In0_c0,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid323_In1_c0,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c0);
   Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid327_In0_c0 <= "" & bh7_w51_2_c0 & bh7_w51_5_c0 & bh7_w51_6_c0 & bh7_w51_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid327_In1_c0 <= "" & bh7_w52_2_c0;
   bh7_w51_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1(0);
   bh7_w52_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1(1);
   bh7_w53_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid327: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid327_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid327_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid329_In0_c0 <= "" & bh7_w52_5_c0 & bh7_w52_6_c0 & bh7_w52_7_c0 & bh7_w52_8_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid329_In1_c0 <= "" & bh7_w53_2_c0;
   bh7_w52_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1(0);
   bh7_w53_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1(1);
   bh7_w54_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid329: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid329_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid329_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid331_In0_c0 <= "" & bh7_w53_5_c0 & bh7_w53_6_c0 & bh7_w53_7_c0 & bh7_w53_8_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid331_In1_c0 <= "" & bh7_w54_2_c0;
   bh7_w53_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1(0);
   bh7_w54_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1(1);
   bh7_w55_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid331: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid331_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid331_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid335_In0_c0 <= "" & bh7_w54_3_c0 & bh7_w54_6_c0 & bh7_w54_7_c0 & bh7_w54_8_c0 & bh7_w54_9_c0 & bh7_w54_10_c0;
   bh7_w54_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1(0);
   bh7_w55_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1(1);
   bh7_w56_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid335: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid335_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid337_In0_c0 <= "" & bh7_w55_2_c0 & bh7_w55_3_c0 & bh7_w55_6_c0 & bh7_w55_7_c0 & bh7_w55_8_c0 & bh7_w55_9_c0;
   bh7_w55_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1(0);
   bh7_w56_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1(1);
   bh7_w57_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid337: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid337_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid339_In0_c0 <= "" & bh7_w56_2_c0 & bh7_w56_5_c0 & bh7_w56_6_c0 & bh7_w56_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid339_In1_c0 <= "" & bh7_w57_2_c0;
   bh7_w56_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1(0);
   bh7_w57_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1(1);
   bh7_w58_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid339: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid339_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid339_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid341_In0_c0 <= "" & bh7_w57_3_c0 & bh7_w57_6_c0 & bh7_w57_7_c0 & bh7_w57_8_c0 & bh7_w57_9_c0 & bh7_w57_10_c0;
   bh7_w57_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1(0);
   bh7_w58_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1(1);
   bh7_w59_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid341: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid341_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid343_In0_c0 <= "" & bh7_w58_1_c0 & bh7_w58_2_c0 & bh7_w58_6_c0 & bh7_w58_7_c0 & bh7_w58_8_c0 & bh7_w58_9_c0;
   bh7_w58_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1(0);
   bh7_w59_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1(1);
   bh7_w60_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid343: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid343_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid345_In0_c0 <= "" & bh7_w59_1_c0 & bh7_w59_5_c0 & bh7_w59_6_c0 & bh7_w59_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid345_In1_c0 <= "" & bh7_w60_1_c0;
   bh7_w59_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1(0);
   bh7_w60_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1(1);
   bh7_w61_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid345: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid345_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid345_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid347_In0_c0 <= "" & bh7_w60_2_c0 & bh7_w60_6_c0 & bh7_w60_7_c0 & bh7_w60_8_c0 & bh7_w60_9_c0 & bh7_w60_10_c0;
   bh7_w60_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1(0);
   bh7_w61_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1(1);
   bh7_w62_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid347: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid347_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid349_In0_c0 <= "" & bh7_w61_1_c0 & bh7_w61_2_c0 & bh7_w61_6_c0 & bh7_w61_7_c0 & bh7_w61_8_c0 & bh7_w61_9_c0;
   bh7_w61_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1(0);
   bh7_w62_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1(1);
   bh7_w63_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid349: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid349_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid351_In0_c0 <= "" & bh7_w62_1_c0 & bh7_w62_5_c0 & bh7_w62_6_c0 & bh7_w62_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid351_In1_c0 <= "" & bh7_w63_1_c0;
   bh7_w62_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1(0);
   bh7_w63_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1(1);
   bh7_w64_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid351: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid351_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid351_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid353_In0_c0 <= "" & bh7_w63_2_c0 & bh7_w63_6_c0 & bh7_w63_7_c0 & bh7_w63_8_c0 & bh7_w63_9_c0 & bh7_w63_10_c0;
   bh7_w63_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1(0);
   bh7_w64_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1(1);
   bh7_w65_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid353: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid353_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid355_In0_c0 <= "" & bh7_w64_1_c0 & bh7_w64_2_c0 & bh7_w64_6_c0 & bh7_w64_7_c0 & bh7_w64_8_c0 & bh7_w64_9_c0;
   bh7_w64_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1(0);
   bh7_w65_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1(1);
   bh7_w66_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid355: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid355_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid357_In0_c0 <= "" & bh7_w65_1_c0 & bh7_w65_4_c0 & bh7_w65_5_c0 & bh7_w65_6_c0 & bh7_w65_7_c0 & bh7_w65_8_c0;
   bh7_w65_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1(0);
   bh7_w66_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1(1);
   bh7_w67_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid357: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid357_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid359_In0_c0 <= "" & bh7_w66_1_c0 & bh7_w66_2_c0 & bh7_w66_5_c0 & bh7_w66_6_c0 & bh7_w66_7_c0 & bh7_w66_8_c0;
   bh7_w66_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1(0);
   bh7_w67_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1(1);
   bh7_w68_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid359: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid359_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid361_In0_c0 <= "" & bh7_w67_1_c0 & bh7_w67_2_c0 & bh7_w67_5_c0 & bh7_w67_6_c0 & bh7_w67_7_c0 & bh7_w67_8_c0;
   bh7_w67_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1(0);
   bh7_w68_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1(1);
   bh7_w69_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid361: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid361_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid363_In0_c0 <= "" & bh7_w68_1_c0 & bh7_w68_4_c0 & bh7_w68_5_c0 & bh7_w68_6_c0 & bh7_w68_7_c0 & bh7_w68_8_c0;
   bh7_w68_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1(0);
   bh7_w69_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1(1);
   bh7_w70_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid363: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid363_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid365_In0_c0 <= "" & bh7_w69_1_c0 & bh7_w69_2_c0 & bh7_w69_5_c0 & bh7_w69_6_c0 & bh7_w69_7_c0 & bh7_w69_8_c0;
   bh7_w69_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1(0);
   bh7_w70_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1(1);
   bh7_w71_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid365: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid365_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid367_In0_c0 <= "" & bh7_w70_1_c0 & bh7_w70_2_c0 & bh7_w70_5_c0 & bh7_w70_6_c0 & bh7_w70_7_c0 & bh7_w70_8_c0;
   bh7_w70_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1(0);
   bh7_w71_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1(1);
   bh7_w72_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid367: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid367_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid369_In0_c0 <= "" & bh7_w71_1_c0 & bh7_w71_4_c0 & bh7_w71_5_c0 & bh7_w71_6_c0 & bh7_w71_7_c0 & bh7_w71_8_c0;
   bh7_w71_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1(0);
   bh7_w72_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1(1);
   bh7_w73_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid369: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid369_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid371_In0_c0 <= "" & bh7_w72_1_c0 & bh7_w72_2_c0 & bh7_w72_5_c0 & bh7_w72_6_c0 & bh7_w72_7_c0 & bh7_w72_8_c0;
   bh7_w72_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1(0);
   bh7_w73_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1(1);
   bh7_w74_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid371: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid371_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid373_In0_c0 <= "" & bh7_w73_1_c0 & bh7_w73_2_c0 & bh7_w73_5_c0 & bh7_w73_6_c0 & bh7_w73_7_c0 & bh7_w73_8_c0;
   bh7_w73_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1(0);
   bh7_w74_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1(1);
   bh7_w75_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid373: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid373_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid375_In0_c0 <= "" & bh7_w74_1_c0 & bh7_w74_4_c0 & bh7_w74_5_c0 & bh7_w74_6_c0 & bh7_w74_7_c0 & bh7_w74_8_c0;
   bh7_w74_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1(0);
   bh7_w75_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1(1);
   bh7_w76_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid375: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid375_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid377_In0_c0 <= "" & bh7_w75_0_c0 & bh7_w75_3_c0 & bh7_w75_4_c0 & bh7_w75_5_c0 & bh7_w75_6_c0 & bh7_w75_7_c0;
   bh7_w75_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1(0);
   bh7_w76_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1(1);
   bh7_w77_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid377: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid377_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid379_In0_c0 <= "" & bh7_w76_0_c0 & bh7_w76_3_c0 & bh7_w76_4_c0 & bh7_w76_5_c0 & bh7_w76_6_c0 & bh7_w76_7_c0;
   bh7_w76_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1(0);
   bh7_w77_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1(1);
   bh7_w78_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid379: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid379_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid381_In0_c0 <= "" & bh7_w77_2_c0 & bh7_w77_3_c0 & bh7_w77_4_c0 & bh7_w77_5_c0 & bh7_w77_6_c0 & bh7_w77_7_c0;
   bh7_w77_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1(0);
   bh7_w78_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1(1);
   bh7_w79_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid381: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid381_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid383_In0_c0 <= "" & bh7_w78_2_c0 & bh7_w78_3_c0 & bh7_w78_4_c0 & bh7_w78_5_c0 & bh7_w78_6_c0 & bh7_w78_7_c0;
   bh7_w78_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1(0);
   bh7_w79_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1(1);
   bh7_w80_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid383: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid383_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid385_In0_c0 <= "" & bh7_w79_2_c0 & bh7_w79_3_c0 & bh7_w79_4_c0 & bh7_w79_5_c0 & bh7_w79_6_c0 & bh7_w79_7_c0;
   bh7_w79_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1(0);
   bh7_w80_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1(1);
   bh7_w81_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid385: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid385_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid387_In0_c0 <= "" & bh7_w80_2_c0 & bh7_w80_3_c0 & bh7_w80_4_c0 & bh7_w80_5_c0 & bh7_w80_6_c0 & bh7_w80_7_c0;
   bh7_w80_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1(0);
   bh7_w81_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1(1);
   bh7_w82_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid387: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid387_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid389_In0_c0 <= "" & bh7_w81_2_c0 & bh7_w81_3_c0 & bh7_w81_4_c0 & bh7_w81_5_c0 & bh7_w81_6_c0 & bh7_w81_7_c0;
   bh7_w81_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1(0);
   bh7_w82_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1(1);
   bh7_w83_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid389: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid389_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid391_In0_c0 <= "" & bh7_w82_1_c0 & bh7_w82_2_c0 & bh7_w82_3_c0 & bh7_w82_4_c0 & bh7_w82_5_c0 & bh7_w82_6_c0;
   bh7_w82_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1(0);
   bh7_w83_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1(1);
   bh7_w84_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid391: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid391_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid393_In0_c0 <= "" & bh7_w83_1_c0 & bh7_w83_2_c0 & bh7_w83_3_c0 & bh7_w83_4_c0 & bh7_w83_5_c0 & bh7_w83_6_c0;
   bh7_w83_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1(0);
   bh7_w84_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1(1);
   bh7_w85_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid393: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid393_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid395_In0_c0 <= "" & bh7_w84_1_c0 & bh7_w84_2_c0 & bh7_w84_3_c0 & bh7_w84_4_c0 & bh7_w84_5_c0 & bh7_w84_6_c0;
   bh7_w84_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1(0);
   bh7_w85_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1(1);
   bh7_w86_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid395: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid395_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid397_In0_c0 <= "" & bh7_w85_1_c0 & bh7_w85_2_c0 & bh7_w85_3_c0 & bh7_w85_4_c0 & bh7_w85_5_c0 & bh7_w85_6_c0;
   bh7_w85_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1(0);
   bh7_w86_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1(1);
   bh7_w87_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid397: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid397_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid401_In0_c0 <= "" & bh7_w86_1_c0 & bh7_w86_2_c0 & bh7_w86_3_c0 & bh7_w86_4_c0 & bh7_w86_5_c0;
   bh7_w86_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1(0);
   bh7_w87_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1(1);
   bh7_w88_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid401: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid401_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid403_In0_c0 <= "" & bh7_w87_1_c0 & bh7_w87_2_c0 & bh7_w87_3_c0 & bh7_w87_4_c0 & bh7_w87_5_c0 & bh7_w87_6_c0;
   bh7_w87_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1(0);
   bh7_w88_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1(1);
   bh7_w89_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid403: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid403_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid405_In0_c0 <= "" & bh7_w88_1_c0 & bh7_w88_2_c0 & bh7_w88_3_c0 & bh7_w88_4_c0 & bh7_w88_5_c0 & bh7_w88_6_c0;
   bh7_w88_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1(0);
   bh7_w89_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1(1);
   bh7_w90_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid405: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid405_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid407_In0_c0 <= "" & bh7_w89_1_c0 & bh7_w89_2_c0 & bh7_w89_3_c0 & bh7_w89_4_c0 & bh7_w89_5_c0;
   bh7_w89_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1(0);
   bh7_w90_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1(1);
   bh7_w91_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid407: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid407_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid409_In0_c0 <= "" & bh7_w90_1_c0 & bh7_w90_2_c0 & bh7_w90_3_c0 & bh7_w90_4_c0 & bh7_w90_5_c0 & bh7_w90_6_c0;
   bh7_w90_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1(0);
   bh7_w91_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1(1);
   bh7_w92_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid409: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid409_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid411_In0_c0 <= "" & bh7_w91_1_c0 & bh7_w91_2_c0 & bh7_w91_3_c0 & bh7_w91_4_c0 & bh7_w91_5_c0 & bh7_w91_6_c0;
   bh7_w91_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1(0);
   bh7_w92_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1(1);
   bh7_w93_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid411: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid411_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid413_In0_c0 <= "" & bh7_w92_1_c0 & bh7_w92_2_c0 & bh7_w92_3_c0 & bh7_w92_4_c0 & bh7_w92_5_c0;
   bh7_w92_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1(0);
   bh7_w93_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1(1);
   bh7_w94_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid413: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid413_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid415_In0_c0 <= "" & bh7_w93_1_c0 & bh7_w93_2_c0 & bh7_w93_3_c0 & bh7_w93_4_c0 & bh7_w93_5_c0 & bh7_w93_6_c0;
   bh7_w93_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1(0);
   bh7_w94_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1(1);
   bh7_w95_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid415: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid415_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid417_In0_c0 <= "" & bh7_w94_1_c0 & bh7_w94_2_c0 & bh7_w94_3_c0 & bh7_w94_4_c0 & bh7_w94_5_c0 & bh7_w94_6_c0;
   bh7_w94_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1(0);
   bh7_w95_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1(1);
   bh7_w96_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid417: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid417_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid419_In0_c0 <= "" & bh7_w95_1_c0 & bh7_w95_2_c0 & bh7_w95_3_c0 & bh7_w95_4_c0 & bh7_w95_5_c0;
   bh7_w95_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1(0);
   bh7_w96_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1(1);
   bh7_w97_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid419: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid419_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid421_In0_c0 <= "" & bh7_w96_1_c0 & bh7_w96_2_c0 & bh7_w96_3_c0 & bh7_w96_4_c0 & bh7_w96_5_c0 & bh7_w96_6_c0;
   bh7_w96_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1(0);
   bh7_w97_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1(1);
   bh7_w98_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid421: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid421_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid423_In0_c0 <= "" & bh7_w97_1_c0 & bh7_w97_2_c0 & bh7_w97_3_c0 & bh7_w97_4_c0 & bh7_w97_5_c0 & bh7_w97_6_c0;
   bh7_w97_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1(0);
   bh7_w98_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1(1);
   bh7_w99_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid423: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid423_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid425_In0_c0 <= "" & bh7_w98_1_c0 & bh7_w98_2_c0 & bh7_w98_3_c0 & bh7_w98_4_c0 & bh7_w98_5_c0;
   bh7_w98_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1(0);
   bh7_w99_7_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1(1);
   bh7_w100_6_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid425: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid425_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid427_In0_c0 <= "" & bh7_w99_0_c0 & bh7_w99_1_c0 & bh7_w99_2_c0 & bh7_w99_3_c0 & bh7_w99_4_c0 & bh7_w99_5_c0;
   bh7_w99_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1(0);
   bh7_w100_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1(1);
   bh7_w101_3_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid427: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid427_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid429_In0_c0 <= "" & bh7_w100_0_c0 & bh7_w100_1_c0 & bh7_w100_2_c0 & bh7_w100_3_c0 & bh7_w100_4_c0 & bh7_w100_5_c0;
   bh7_w100_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1(0);
   bh7_w101_4_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1(1);
   bh7_w102_4_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid429: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid429_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid433_In0_c0 <= "" & bh7_w101_0_c0 & bh7_w101_1_c0 & bh7_w101_2_c0;
   bh7_w101_5_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1(0);
   bh7_w102_5_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid433: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid433_In0_c0,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c0);
   Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid435_In0_c0 <= "" & bh7_w102_0_c0 & bh7_w102_1_c0 & bh7_w102_2_c0 & bh7_w102_3_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid435_In1_c0 <= "" & bh7_w103_0_c0;
   bh7_w102_6_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1(0);
   bh7_w103_2_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1(1);
   bh7_w104_1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid435: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid435_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid435_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid437_In0_c1 <= "" & bh7_w51_9_c1 & bh7_w51_8_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid437_In1_c1 <= "" & bh7_w52_10_c1 & bh7_w52_9_c1;
   bh7_w51_10_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1(0);
   bh7_w52_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1(1);
   bh7_w53_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid437: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid437_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid437_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_copy438_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_copy438_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid439_In0_c1 <= "" & bh7_w53_11_c1 & bh7_w53_10_c1 & bh7_w53_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid439_In1_c1 <= "" & bh7_w54_12_c1 & bh7_w54_11_c1;
   bh7_w53_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1(0);
   bh7_w54_14_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1(1);
   bh7_w55_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid439: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid439_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid439_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_copy440_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_copy440_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid441_In0_c1 <= "" & bh7_w55_10_c1 & bh7_w55_12_c1 & bh7_w55_11_c1;
   bh7_w55_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1(0);
   bh7_w56_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid441: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid441_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_copy442_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_copy442_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid443_In0_c1 <= "" & bh7_w56_8_c1 & bh7_w56_11_c1 & bh7_w56_10_c1 & bh7_w56_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c0 <= "" & "0";
   bh7_w56_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1(0);
   bh7_w57_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1(1);
   bh7_w58_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid443: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid443_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_copy444_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_copy444_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid445_In0_c1 <= "" & bh7_w57_12_c1 & bh7_w57_13_c1 & bh7_w57_11_c1;
   bh7_w57_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1(0);
   bh7_w58_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid445: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid445_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_copy446_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_copy446_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid447_In0_c1 <= "" & bh7_w58_10_c1 & bh7_w58_12_c1 & bh7_w58_11_c1;
   bh7_w58_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1(0);
   bh7_w59_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid447: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid447_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_copy448_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_copy448_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid449_In0_c1 <= "" & bh7_w59_8_c1 & bh7_w59_11_c1 & bh7_w59_10_c1 & bh7_w59_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c0 <= "" & "0";
   bh7_w59_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1(0);
   bh7_w60_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1(1);
   bh7_w61_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid449: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid449_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_copy450_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_copy450_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid451_In0_c1 <= "" & bh7_w60_12_c1 & bh7_w60_13_c1 & bh7_w60_11_c1;
   bh7_w60_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1(0);
   bh7_w61_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid451: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid451_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_copy452_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_copy452_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid453_In0_c1 <= "" & bh7_w61_10_c1 & bh7_w61_12_c1 & bh7_w61_11_c1;
   bh7_w61_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1(0);
   bh7_w62_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid453: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid453_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_copy454_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_copy454_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid455_In0_c1 <= "" & bh7_w62_8_c1 & bh7_w62_11_c1 & bh7_w62_10_c1 & bh7_w62_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c0 <= "" & "0";
   bh7_w62_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1(0);
   bh7_w63_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1(1);
   bh7_w64_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid455: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid455_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_copy456_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_copy456_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid457_In0_c1 <= "" & bh7_w63_12_c1 & bh7_w63_13_c1 & bh7_w63_11_c1;
   bh7_w63_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1(0);
   bh7_w64_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid457: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid457_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_copy458_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_copy458_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid459_In0_c1 <= "" & bh7_w64_10_c1 & bh7_w64_12_c1 & bh7_w64_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid459_In1_c1 <= "" & bh7_w65_11_c1 & bh7_w65_10_c1;
   bh7_w64_15_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1(0);
   bh7_w65_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1(1);
   bh7_w66_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid459: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid459_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid459_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_copy460_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_copy460_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid461_In0_c1 <= "" & bh7_w66_9_c1 & bh7_w66_12_c1 & bh7_w66_11_c1 & bh7_w66_10_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c0 <= "" & "0";
   bh7_w66_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1(0);
   bh7_w67_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1(1);
   bh7_w68_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid461: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid461_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_copy462_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_copy462_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid463_In0_c1 <= "" & bh7_w67_11_c1 & bh7_w67_10_c1 & bh7_w67_9_c1;
   bh7_w67_13_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1(0);
   bh7_w68_13_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid463: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid463_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_copy464_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_copy464_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid465_In0_c1 <= "" & bh7_w68_11_c1 & bh7_w68_10_c1 & bh7_w68_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid465_In1_c1 <= "" & bh7_w69_11_c1 & bh7_w69_10_c1;
   bh7_w68_14_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1(0);
   bh7_w69_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1(1);
   bh7_w70_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid465: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid465_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid465_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_copy466_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_copy466_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid467_In0_c1 <= "" & bh7_w70_11_c1 & bh7_w70_10_c1 & bh7_w70_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid467_In1_c1 <= "" & bh7_w71_11_c1 & bh7_w71_10_c1;
   bh7_w70_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1(0);
   bh7_w71_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1(1);
   bh7_w72_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid467: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid467_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid467_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_copy468_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_copy468_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid469_In0_c1 <= "" & bh7_w72_11_c1 & bh7_w72_10_c1 & bh7_w72_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid469_In1_c1 <= "" & bh7_w73_11_c1 & bh7_w73_10_c1;
   bh7_w72_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1(0);
   bh7_w73_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1(1);
   bh7_w74_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid469: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid469_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid469_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_copy470_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_copy470_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid471_In0_c1 <= "" & bh7_w74_11_c1 & bh7_w74_10_c1 & bh7_w74_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid471_In1_c1 <= "" & bh7_w75_10_c1 & bh7_w75_9_c1;
   bh7_w74_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1(0);
   bh7_w75_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1(1);
   bh7_w76_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid471: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid471_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid471_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_copy472_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_copy472_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid473_In0_c1 <= "" & bh7_w76_10_c1 & bh7_w76_9_c1 & bh7_w76_8_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid473_In1_c1 <= "" & bh7_w77_10_c1 & bh7_w77_9_c1;
   bh7_w76_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1(0);
   bh7_w77_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1(1);
   bh7_w78_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid473: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid473_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid473_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_copy474_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_copy474_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid475_In0_c1 <= "" & bh7_w78_10_c1 & bh7_w78_9_c1 & bh7_w78_8_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid475_In1_c1 <= "" & bh7_w79_10_c1 & bh7_w79_9_c1;
   bh7_w78_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1(0);
   bh7_w79_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1(1);
   bh7_w80_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid475: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid475_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid475_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_copy476_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_copy476_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid477_In0_c1 <= "" & bh7_w80_10_c1 & bh7_w80_9_c1 & bh7_w80_8_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid477_In1_c1 <= "" & bh7_w81_10_c1 & bh7_w81_9_c1;
   bh7_w80_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1(0);
   bh7_w81_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1(1);
   bh7_w82_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid477: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid477_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid477_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_copy478_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_copy478_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid479_In0_c1 <= "" & bh7_w82_7_c1 & bh7_w82_10_c1 & bh7_w82_9_c1 & bh7_w82_8_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c0 <= "" & "0";
   bh7_w82_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1(0);
   bh7_w83_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1(1);
   bh7_w84_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid479: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid479_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_copy480_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_copy480_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid481_In0_c1 <= "" & bh7_w83_9_c1 & bh7_w83_8_c1 & bh7_w83_7_c1;
   bh7_w83_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1(0);
   bh7_w84_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid481: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid481_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_copy482_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_copy482_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid483_In0_c1 <= "" & bh7_w84_9_c1 & bh7_w84_8_c1 & bh7_w84_7_c1;
   bh7_w84_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1(0);
   bh7_w85_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid483: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid483_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_copy484_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_copy484_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid485_In0_c1 <= "" & bh7_w85_7_c1 & bh7_w85_10_c1 & bh7_w85_9_c1 & bh7_w85_8_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c0 <= "" & "0";
   bh7_w85_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1(0);
   bh7_w86_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1(1);
   bh7_w87_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid485: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid485_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_copy486_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_copy486_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid487_In0_c1 <= "" & bh7_w86_8_c1 & bh7_w86_7_c1 & bh7_w86_6_c1;
   bh7_w86_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1(0);
   bh7_w87_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid487: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid487_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_copy488_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_copy488_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid489_In0_c1 <= "" & bh7_w87_8_c1 & bh7_w87_9_c1 & bh7_w87_7_c1;
   bh7_w87_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1(0);
   bh7_w88_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid489: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid489_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_copy490_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_copy490_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid491_In0_c1 <= "" & bh7_w88_7_c1 & bh7_w88_8_c1 & bh7_w88_10_c1 & bh7_w88_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c0 <= "" & "0";
   bh7_w88_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1(0);
   bh7_w89_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1(1);
   bh7_w90_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid491: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid491_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_copy492_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_copy492_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid493_In0_c1 <= "" & bh7_w89_8_c1 & bh7_w89_7_c1 & bh7_w89_6_c1;
   bh7_w89_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1(0);
   bh7_w90_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid493: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid493_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_copy494_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_copy494_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid495_In0_c1 <= "" & bh7_w90_8_c1 & bh7_w90_9_c1 & bh7_w90_7_c1;
   bh7_w90_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1(0);
   bh7_w91_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid495: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid495_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_copy496_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_copy496_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid497_In0_c1 <= "" & bh7_w91_7_c1 & bh7_w91_8_c1 & bh7_w91_10_c1 & bh7_w91_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c0 <= "" & "0";
   bh7_w91_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1(0);
   bh7_w92_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1(1);
   bh7_w93_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid497: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid497_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_copy498_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_copy498_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid499_In0_c1 <= "" & bh7_w92_8_c1 & bh7_w92_7_c1 & bh7_w92_6_c1;
   bh7_w92_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1(0);
   bh7_w93_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid499: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid499_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_copy500_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_copy500_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid501_In0_c1 <= "" & bh7_w93_8_c1 & bh7_w93_9_c1 & bh7_w93_7_c1;
   bh7_w93_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1(0);
   bh7_w94_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid501: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid501_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_copy502_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_copy502_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid503_In0_c1 <= "" & bh7_w94_7_c1 & bh7_w94_8_c1 & bh7_w94_10_c1 & bh7_w94_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c0 <= "" & "0";
   bh7_w94_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1(0);
   bh7_w95_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1(1);
   bh7_w96_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid503: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid503_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_copy504_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_copy504_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid505_In0_c1 <= "" & bh7_w95_8_c1 & bh7_w95_7_c1 & bh7_w95_6_c1;
   bh7_w95_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1(0);
   bh7_w96_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid505: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid505_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_copy506_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_copy506_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid507_In0_c1 <= "" & bh7_w96_8_c1 & bh7_w96_9_c1 & bh7_w96_7_c1;
   bh7_w96_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1(0);
   bh7_w97_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid507: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid507_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_copy508_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_copy508_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid509_In0_c1 <= "" & bh7_w97_7_c1 & bh7_w97_8_c1 & bh7_w97_10_c1 & bh7_w97_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c0 <= "" & "0";
   bh7_w97_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1(0);
   bh7_w98_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1(1);
   bh7_w99_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid509: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid509_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_copy510_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_copy510_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid511_In0_c1 <= "" & bh7_w98_8_c1 & bh7_w98_7_c1 & bh7_w98_6_c1;
   bh7_w98_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1(0);
   bh7_w99_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid511: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid511_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_copy512_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_copy512_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid513_In0_c1 <= "" & bh7_w99_7_c1 & bh7_w99_8_c1 & bh7_w99_6_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid513_In1_c1 <= "" & bh7_w100_6_c1 & bh7_w100_8_c1;
   bh7_w99_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1(0);
   bh7_w100_9_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1(1);
   bh7_w101_6_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid513: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid513_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid513_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_copy514_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_copy514_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid515_In0_c1 <= "" & bh7_w101_5_c1 & bh7_w101_4_c1 & bh7_w101_3_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid515_In1_c1 <= "" & bh7_w102_6_c1 & bh7_w102_5_c1;
   bh7_w101_7_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1(0);
   bh7_w102_7_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1(1);
   bh7_w103_3_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid515: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid515_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid515_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_copy516_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_copy516_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid517_In0_c1 <= "" & bh7_w103_1_c1 & bh7_w103_2_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid517_In1_c1 <= "" & bh7_w104_0_c1 & bh7_w104_1_c1;
   bh7_w103_4_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1(0);
   bh7_w104_2_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1(1);
   bh7_w105_1_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid517: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid517_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid517_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_copy518_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_copy518_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid519_In0_c1 <= "" & bh7_w53_13_c1 & bh7_w53_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid519_In1_c1 <= "" & bh7_w54_13_c1 & bh7_w54_14_c1;
   bh7_w53_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2(0);
   bh7_w54_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2(1);
   bh7_w55_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid519: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid519_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid519_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid521_In0_c1 <= "" & bh7_w55_13_c1 & bh7_w55_14_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid521_In1_c1 <= "" & bh7_w56_13_c1 & bh7_w56_12_c1;
   bh7_w55_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2(0);
   bh7_w56_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2(1);
   bh7_w57_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid521: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid521_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid521_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid523_In0_c1 <= "" & bh7_w57_14_c1 & bh7_w57_15_c1 & "0";
   bh7_w57_17_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2(0);
   bh7_w58_16_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid523: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid523_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid525_In0_c1 <= "" & bh7_w58_13_c1 & bh7_w58_15_c1 & bh7_w58_14_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid525_In1_c1 <= "" & bh7_w59_13_c1 & bh7_w59_12_c1;
   bh7_w58_17_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2(0);
   bh7_w59_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2(1);
   bh7_w60_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid525: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid525_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid525_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid527_In0_c1 <= "" & bh7_w60_14_c1 & bh7_w60_15_c1 & "0";
   bh7_w60_17_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2(0);
   bh7_w61_16_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid527: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid527_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid529_In0_c1 <= "" & bh7_w61_13_c1 & bh7_w61_15_c1 & bh7_w61_14_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid529_In1_c1 <= "" & bh7_w62_13_c1 & bh7_w62_12_c1;
   bh7_w61_17_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2(0);
   bh7_w62_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2(1);
   bh7_w63_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid529: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid529_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid529_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid531_In0_c1 <= "" & bh7_w63_14_c1 & bh7_w63_15_c1 & "0";
   bh7_w63_17_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2(0);
   bh7_w64_16_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid531: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid531_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid533_In0_c1 <= "" & bh7_w64_13_c1 & bh7_w64_15_c1 & bh7_w64_14_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid533_In1_c1 <= "" & bh7_w65_9_c1 & bh7_w65_12_c1;
   bh7_w64_17_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2(0);
   bh7_w65_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2(1);
   bh7_w66_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid533: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid533_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid533_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid535_In0_c1 <= "" & bh7_w66_14_c1 & bh7_w66_13_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid535_In1_c1 <= "" & bh7_w67_12_c1 & bh7_w67_13_c1;
   bh7_w66_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2(0);
   bh7_w67_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2(1);
   bh7_w68_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid535: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid535_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid535_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid537_In0_c1 <= "" & bh7_w68_12_c1 & bh7_w68_14_c1 & bh7_w68_13_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid537_In1_c1 <= "" & bh7_w69_9_c1 & bh7_w69_12_c1;
   bh7_w68_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2(0);
   bh7_w69_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2(1);
   bh7_w70_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid537: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid537_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid537_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid539_In0_c1 <= "" & bh7_w70_13_c1 & bh7_w70_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid539_In1_c1 <= "" & bh7_w71_9_c1 & bh7_w71_12_c1;
   bh7_w70_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2(0);
   bh7_w71_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2(1);
   bh7_w72_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid539: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid539_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid539_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid541_In0_c1 <= "" & bh7_w72_13_c1 & bh7_w72_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid541_In1_c1 <= "" & bh7_w73_9_c1 & bh7_w73_12_c1;
   bh7_w72_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2(0);
   bh7_w73_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2(1);
   bh7_w74_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid541: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid541_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid541_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid543_In0_c1 <= "" & bh7_w74_13_c1 & bh7_w74_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid543_In1_c1 <= "" & bh7_w75_8_c1 & bh7_w75_11_c1;
   bh7_w74_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2(0);
   bh7_w75_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2(1);
   bh7_w76_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid543: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid543_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid543_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid545_In0_c1 <= "" & bh7_w76_12_c1 & bh7_w76_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid545_In1_c1 <= "" & bh7_w77_8_c1 & bh7_w77_11_c1;
   bh7_w76_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2(0);
   bh7_w77_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2(1);
   bh7_w78_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid545: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid545_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid545_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid547_In0_c1 <= "" & bh7_w78_12_c1 & bh7_w78_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid547_In1_c1 <= "" & bh7_w79_8_c1 & bh7_w79_11_c1;
   bh7_w78_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2(0);
   bh7_w79_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2(1);
   bh7_w80_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid547: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid547_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid547_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid549_In0_c1 <= "" & bh7_w80_12_c1 & bh7_w80_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid549_In1_c1 <= "" & bh7_w81_8_c1 & bh7_w81_11_c1;
   bh7_w80_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2(0);
   bh7_w81_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2(1);
   bh7_w82_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid549: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid549_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid549_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid551_In0_c1 <= "" & bh7_w82_12_c1 & bh7_w82_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid551_In1_c1 <= "" & bh7_w83_10_c1 & bh7_w83_11_c1;
   bh7_w82_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2(0);
   bh7_w83_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2(1);
   bh7_w84_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid551: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid551_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid551_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid553_In0_c1 <= "" & bh7_w84_10_c1 & bh7_w84_12_c1 & bh7_w84_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid553_In1_c1 <= "" & bh7_w85_12_c1 & bh7_w85_11_c1;
   bh7_w84_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2(0);
   bh7_w85_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2(1);
   bh7_w86_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid553: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid553_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid553_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid555_In0_c1 <= "" & bh7_w86_9_c1 & bh7_w86_10_c1 & "0";
   bh7_w86_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2(0);
   bh7_w87_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid555: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid555_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid557_In0_c1 <= "" & bh7_w87_10_c1 & bh7_w87_12_c1 & bh7_w87_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid557_In1_c1 <= "" & bh7_w88_12_c1 & bh7_w88_11_c1;
   bh7_w87_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2(0);
   bh7_w88_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2(1);
   bh7_w89_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid557: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid557_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid557_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid559_In0_c1 <= "" & bh7_w89_9_c1 & bh7_w89_10_c1 & "0";
   bh7_w89_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2(0);
   bh7_w90_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid559: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid559_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid561_In0_c1 <= "" & bh7_w90_10_c1 & bh7_w90_12_c1 & bh7_w90_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid561_In1_c1 <= "" & bh7_w91_12_c1 & bh7_w91_11_c1;
   bh7_w90_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2(0);
   bh7_w91_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2(1);
   bh7_w92_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid561: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid561_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid561_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid563_In0_c1 <= "" & bh7_w92_9_c1 & bh7_w92_10_c1 & "0";
   bh7_w92_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2(0);
   bh7_w93_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid563: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid563_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid565_In0_c1 <= "" & bh7_w93_10_c1 & bh7_w93_12_c1 & bh7_w93_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid565_In1_c1 <= "" & bh7_w94_12_c1 & bh7_w94_11_c1;
   bh7_w93_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2(0);
   bh7_w94_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2(1);
   bh7_w95_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid565: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid565_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid565_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid567_In0_c1 <= "" & bh7_w95_9_c1 & bh7_w95_10_c1 & "0";
   bh7_w95_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2(0);
   bh7_w96_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid567: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid567_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid569_In0_c1 <= "" & bh7_w96_10_c1 & bh7_w96_12_c1 & bh7_w96_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid569_In1_c1 <= "" & bh7_w97_12_c1 & bh7_w97_11_c1;
   bh7_w96_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2(0);
   bh7_w97_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2(1);
   bh7_w98_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid569: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid569_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid569_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid571_In0_c1 <= "" & bh7_w98_9_c1 & bh7_w98_10_c1 & "0";
   bh7_w98_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2(0);
   bh7_w99_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid571: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid571_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid573_In0_c1 <= "" & bh7_w99_9_c1 & bh7_w99_11_c1 & bh7_w99_10_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid573_In1_c1 <= "" & bh7_w100_7_c1 & bh7_w100_9_c1;
   bh7_w99_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2(0);
   bh7_w100_10_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2(1);
   bh7_w101_8_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid573: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid573_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid573_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid575_In0_c1 <= "" & bh7_w101_7_c1 & bh7_w101_6_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid575_In1_c1 <= "" & bh7_w102_4_c1 & bh7_w102_7_c1;
   bh7_w101_9_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2(0);
   bh7_w102_8_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2(1);
   bh7_w103_5_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid575: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid575_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid575_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid577_In0_c1 <= "" & bh7_w103_4_c1 & bh7_w103_3_c1 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid577_In1_c1 <= "" & bh7_w104_2_c1;
   bh7_w103_6_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2(0);
   bh7_w104_3_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2(1);
   bh7_w105_2_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid577: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid577_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid577_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid579_In0_c1 <= "" & bh7_w105_0_c1 & bh7_w105_1_c1 & "0";
   bh7_w105_3_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_c2(0);
   Compressor_3_2_Freq800_uid432_uid579: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid579_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid581_In0_c2 <= "" & bh7_w55_16_c2 & bh7_w55_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid581_In1_c2 <= "" & bh7_w56_14_c2;
   bh7_w55_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2(0);
   bh7_w56_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2(1);
   bh7_w57_18_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid581: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid581_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid581_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_copy582_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_copy582_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid583_In0_c2 <= "" & bh7_w57_16_c2 & bh7_w57_17_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid583_In1_c2 <= "" & bh7_w58_16_c2 & bh7_w58_17_c2;
   bh7_w57_19_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2(0);
   bh7_w58_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2(1);
   bh7_w59_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid583: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid583_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid583_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_copy584_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_copy584_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid585_In0_c2 <= "" & bh7_w60_16_c2 & bh7_w60_17_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid585_In1_c2 <= "" & bh7_w61_16_c2 & bh7_w61_17_c2;
   bh7_w60_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2(0);
   bh7_w61_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2(1);
   bh7_w62_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid585: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid585_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid585_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_copy586_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_copy586_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid587_In0_c2 <= "" & bh7_w63_16_c2 & bh7_w63_17_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid587_In1_c2 <= "" & bh7_w64_16_c2 & bh7_w64_17_c2;
   bh7_w63_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2(0);
   bh7_w64_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2(1);
   bh7_w65_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid587: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid587_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid587_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_copy588_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_copy588_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid589_In0_c2 <= "" & bh7_w66_15_c2 & bh7_w66_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid589_In1_c2 <= "" & bh7_w67_14_c2;
   bh7_w66_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2(0);
   bh7_w67_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2(1);
   bh7_w68_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid589: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid589_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid589_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_copy590_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_copy590_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid591_In0_c2 <= "" & bh7_w68_15_c2 & bh7_w68_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid591_In1_c2 <= "" & bh7_w69_13_c2;
   bh7_w68_18_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2(0);
   bh7_w69_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2(1);
   bh7_w70_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid591: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid591_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid591_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_copy592_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_copy592_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid593_In0_c2 <= "" & bh7_w70_14_c2 & bh7_w70_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid593_In1_c2 <= "" & bh7_w71_13_c2;
   bh7_w70_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2(0);
   bh7_w71_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2(1);
   bh7_w72_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid593: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid593_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid593_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_copy594_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_copy594_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid595_In0_c2 <= "" & bh7_w72_15_c2 & bh7_w72_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid595_In1_c2 <= "" & bh7_w73_13_c2;
   bh7_w72_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2(0);
   bh7_w73_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2(1);
   bh7_w74_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid595: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid595_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid595_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_copy596_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_copy596_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid597_In0_c2 <= "" & bh7_w74_15_c2 & bh7_w74_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid597_In1_c2 <= "" & bh7_w75_12_c2;
   bh7_w74_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2(0);
   bh7_w75_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2(1);
   bh7_w76_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid597: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid597_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid597_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_copy598_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_copy598_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid599_In0_c2 <= "" & bh7_w76_14_c2 & bh7_w76_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid599_In1_c2 <= "" & bh7_w77_12_c2;
   bh7_w76_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2(0);
   bh7_w77_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2(1);
   bh7_w78_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid599: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid599_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid599_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_copy600_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_copy600_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid601_In0_c2 <= "" & bh7_w78_14_c2 & bh7_w78_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid601_In1_c2 <= "" & bh7_w79_12_c2;
   bh7_w78_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2(0);
   bh7_w79_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2(1);
   bh7_w80_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid601: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid601_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid601_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_copy602_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_copy602_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid603_In0_c2 <= "" & bh7_w80_14_c2 & bh7_w80_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid603_In1_c2 <= "" & bh7_w81_12_c2;
   bh7_w80_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2(0);
   bh7_w81_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2(1);
   bh7_w82_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid603: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid603_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid603_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_copy604_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_copy604_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid605_In0_c2 <= "" & bh7_w82_14_c2 & bh7_w82_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid605_In1_c2 <= "" & bh7_w83_12_c2;
   bh7_w82_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2(0);
   bh7_w83_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2(1);
   bh7_w84_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid605: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid605_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid605_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_copy606_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_copy606_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid607_In0_c2 <= "" & bh7_w84_13_c2 & bh7_w84_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid607_In1_c2 <= "" & bh7_w85_13_c2;
   bh7_w84_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2(0);
   bh7_w85_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2(1);
   bh7_w86_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid607: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid607_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid607_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_copy608_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_copy608_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid609_In0_c2 <= "" & bh7_w86_11_c2 & bh7_w86_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid609_In1_c2 <= "" & bh7_w87_13_c2 & bh7_w87_14_c2;
   bh7_w86_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2(0);
   bh7_w87_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2(1);
   bh7_w88_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid609: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid609_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid609_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_copy610_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_copy610_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid611_In0_c2 <= "" & bh7_w89_11_c2 & bh7_w89_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid611_In1_c2 <= "" & bh7_w90_13_c2 & bh7_w90_14_c2;
   bh7_w89_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2(0);
   bh7_w90_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2(1);
   bh7_w91_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid611: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid611_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid611_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_copy612_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_copy612_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid613_In0_c2 <= "" & bh7_w92_11_c2 & bh7_w92_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid613_In1_c2 <= "" & bh7_w93_13_c2 & bh7_w93_14_c2;
   bh7_w92_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2(0);
   bh7_w93_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2(1);
   bh7_w94_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid613: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid613_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid613_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_copy614_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_copy614_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid615_In0_c2 <= "" & bh7_w95_11_c2 & bh7_w95_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid615_In1_c2 <= "" & bh7_w96_13_c2 & bh7_w96_14_c2;
   bh7_w95_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2(0);
   bh7_w96_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2(1);
   bh7_w97_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid615: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid615_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid615_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_copy616_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_copy616_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid617_In0_c2 <= "" & bh7_w98_11_c2 & bh7_w98_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid617_In1_c2 <= "" & bh7_w99_12_c2 & bh7_w99_13_c2;
   bh7_w98_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2(0);
   bh7_w99_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2(1);
   bh7_w100_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid617: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid617_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid617_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_copy618_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_copy618_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid619_In0_c2 <= "" & bh7_w101_8_c2 & bh7_w101_9_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid619_In1_c2 <= "" & bh7_w102_8_c2;
   bh7_w101_10_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2(0);
   bh7_w102_9_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2(1);
   bh7_w103_7_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid619: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid619_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid619_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_copy620_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_copy620_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid621_In0_c2 <= "" & bh7_w103_6_c2 & bh7_w103_5_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid621_In1_c2 <= "" & bh7_w104_3_c2;
   bh7_w103_8_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2(0);
   bh7_w104_4_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2(1);
   bh7_w105_4_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid621: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid621_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid621_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_copy622_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_copy622_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid623_In0_c2 <= "" & bh7_w105_3_c2 & bh7_w105_2_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c0 <= "" & "0";
   bh7_w105_5_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_c2(0);
   Compressor_14_3_Freq800_uid326_uid623: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid623_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_copy624_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_copy624_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid625_In0_c2 <= "" & bh7_w57_18_c2 & bh7_w57_19_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid625_In1_c2 <= "" & bh7_w58_18_c2;
   bh7_w57_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3(0);
   bh7_w58_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3(1);
   bh7_w59_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid625: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid625_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid625_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid627_In0_c2 <= "" & bh7_w59_14_c2 & bh7_w59_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid627_In1_c2 <= "" & bh7_w60_18_c2;
   bh7_w59_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3(0);
   bh7_w60_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3(1);
   bh7_w61_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid627: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid627_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid627_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid629_In0_c2 <= "" & bh7_w62_14_c2 & bh7_w62_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid629_In1_c2 <= "" & bh7_w63_18_c2;
   bh7_w62_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3(0);
   bh7_w63_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3(1);
   bh7_w64_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid629: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid629_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid629_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid631_In0_c2 <= "" & bh7_w65_13_c2 & bh7_w65_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid631_In1_c2 <= "" & bh7_w66_17_c2;
   bh7_w65_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3(0);
   bh7_w66_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3(1);
   bh7_w67_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid631: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid631_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid631_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid633_In0_c2 <= "" & bh7_w68_17_c2 & bh7_w68_18_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid633_In1_c2 <= "" & bh7_w69_14_c2;
   bh7_w68_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3(0);
   bh7_w69_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3(1);
   bh7_w70_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid633: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid633_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid633_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid635_In0_c2 <= "" & bh7_w70_16_c2 & bh7_w70_17_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid635_In1_c2 <= "" & bh7_w71_14_c2;
   bh7_w70_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3(0);
   bh7_w71_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3(1);
   bh7_w72_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid635: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid635_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid635_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid637_In0_c2 <= "" & bh7_w72_16_c2 & bh7_w72_17_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid637_In1_c2 <= "" & bh7_w73_14_c2;
   bh7_w72_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3(0);
   bh7_w73_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3(1);
   bh7_w74_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid637: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid637_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid637_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid639_In0_c2 <= "" & bh7_w74_17_c2 & bh7_w74_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid639_In1_c2 <= "" & bh7_w75_13_c2;
   bh7_w74_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3(0);
   bh7_w75_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3(1);
   bh7_w76_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid639: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid639_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid639_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid641_In0_c2 <= "" & bh7_w76_16_c2 & bh7_w76_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid641_In1_c2 <= "" & bh7_w77_13_c2;
   bh7_w76_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3(0);
   bh7_w77_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3(1);
   bh7_w78_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid641: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid641_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid641_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid643_In0_c2 <= "" & bh7_w78_16_c2 & bh7_w78_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid643_In1_c2 <= "" & bh7_w79_13_c2;
   bh7_w78_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3(0);
   bh7_w79_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3(1);
   bh7_w80_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid643: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid643_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid643_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid645_In0_c2 <= "" & bh7_w80_16_c2 & bh7_w80_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid645_In1_c2 <= "" & bh7_w81_13_c2;
   bh7_w80_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3(0);
   bh7_w81_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3(1);
   bh7_w82_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid645: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid645_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid645_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid647_In0_c2 <= "" & bh7_w82_16_c2 & bh7_w82_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid647_In1_c2 <= "" & bh7_w83_13_c2;
   bh7_w82_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3(0);
   bh7_w83_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3(1);
   bh7_w84_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid647: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid647_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid647_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid649_In0_c2 <= "" & bh7_w84_15_c2 & bh7_w84_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid649_In1_c2 <= "" & bh7_w85_14_c2;
   bh7_w84_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3(0);
   bh7_w85_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3(1);
   bh7_w86_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid649: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid649_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid649_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid651_In0_c2 <= "" & bh7_w86_13_c2 & bh7_w86_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid651_In1_c2 <= "" & bh7_w87_15_c2;
   bh7_w86_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3(0);
   bh7_w87_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3(1);
   bh7_w88_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid651: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid651_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid651_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid653_In0_c2 <= "" & bh7_w88_13_c2 & bh7_w88_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid653_In1_c2 <= "" & bh7_w89_13_c2;
   bh7_w88_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3(0);
   bh7_w89_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3(1);
   bh7_w90_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid653: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid653_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid653_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid655_In0_c2 <= "" & bh7_w91_13_c2 & bh7_w91_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid655_In1_c2 <= "" & bh7_w92_13_c2;
   bh7_w91_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3(0);
   bh7_w92_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3(1);
   bh7_w93_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid655: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid655_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid655_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid657_In0_c2 <= "" & bh7_w94_13_c2 & bh7_w94_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid657_In1_c2 <= "" & bh7_w95_13_c2;
   bh7_w94_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3(0);
   bh7_w95_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3(1);
   bh7_w96_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid657: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid657_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid657_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid659_In0_c2 <= "" & bh7_w97_13_c2 & bh7_w97_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid659_In1_c2 <= "" & bh7_w98_13_c2;
   bh7_w97_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3(0);
   bh7_w98_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3(1);
   bh7_w99_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid659: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid659_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid659_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid661_In0_c2 <= "" & bh7_w100_10_c2 & bh7_w100_11_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid661_In1_c2 <= "" & bh7_w101_10_c2;
   bh7_w100_12_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3(0);
   bh7_w101_11_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3(1);
   bh7_w102_10_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid661: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid661_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid661_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid663_In0_c2 <= "" & bh7_w103_7_c2 & bh7_w103_8_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid663_In1_c2 <= "" & bh7_w104_4_c2;
   bh7_w103_9_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3(0);
   bh7_w104_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3(1);
   bh7_w105_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid663: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid663_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid663_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid665_In0_c2 <= "" & bh7_w105_5_c2 & bh7_w105_4_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c0 <= "" & "0";
   bh7_w105_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_c3(0);
   Compressor_14_3_Freq800_uid326_uid665: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid665_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid667_In0_c2 <= "" & bh7_w17_0_c2 & bh7_w17_1_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid667_In1_c2 <= "" & bh7_w18_0_c2 & bh7_w18_1_c2;
   bh7_w17_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3(0);
   bh7_w18_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3(1);
   bh7_w19_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid667: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid667_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid667_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid669_In0_c2 <= "" & bh7_w19_0_c2 & bh7_w19_1_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid669_In1_c2 <= "" & bh7_w20_0_c2 & bh7_w20_1_c2;
   bh7_w19_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3(0);
   bh7_w20_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3(1);
   bh7_w21_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid669: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid669_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid669_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid671_In0_c2 <= "" & bh7_w21_0_c2 & bh7_w21_1_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid671_In1_c2 <= "" & bh7_w22_0_c2 & bh7_w22_1_c2;
   bh7_w21_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3(0);
   bh7_w22_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3(1);
   bh7_w23_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid671: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid671_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid671_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid673_In0_c2 <= "" & bh7_w23_0_c2 & bh7_w23_1_c2 & "0";
   bh7_w23_3_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3(0);
   bh7_w24_3_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid673: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid673_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid675_In0_c2 <= "" & bh7_w24_0_c2 & bh7_w24_1_c2 & bh7_w24_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid675_In1_c2 <= "" & bh7_w25_0_c2 & bh7_w25_1_c2;
   bh7_w24_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3(0);
   bh7_w25_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3(1);
   bh7_w26_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid675: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid675_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid675_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid677_In0_c2 <= "" & bh7_w26_0_c2 & bh7_w26_1_c2 & bh7_w26_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid677_In1_c2 <= "" & bh7_w27_0_c2 & bh7_w27_1_c2;
   bh7_w26_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3(0);
   bh7_w27_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3(1);
   bh7_w28_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid677: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid677_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid677_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid679_In0_c2 <= "" & bh7_w28_0_c2 & bh7_w28_1_c2 & bh7_w28_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid679_In1_c2 <= "" & bh7_w29_0_c2 & bh7_w29_1_c2;
   bh7_w28_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3(0);
   bh7_w29_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3(1);
   bh7_w30_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid679: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid679_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid679_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid681_In0_c2 <= "" & bh7_w30_0_c2 & bh7_w30_1_c2 & bh7_w30_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid681_In1_c2 <= "" & bh7_w31_0_c2 & bh7_w31_1_c2;
   bh7_w30_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3(0);
   bh7_w31_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3(1);
   bh7_w32_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid681: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid681_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid681_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid683_In0_c2 <= "" & bh7_w32_0_c2 & bh7_w32_1_c2 & bh7_w32_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid683_In1_c2 <= "" & bh7_w33_0_c2 & bh7_w33_1_c2;
   bh7_w32_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3(0);
   bh7_w33_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3(1);
   bh7_w34_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid683: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid683_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid683_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid685_In0_c2 <= "" & bh7_w34_0_c2 & bh7_w34_1_c2 & bh7_w34_2_c2 & bh7_w34_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid685_In1_c2 <= "" & bh7_w35_0_c2;
   bh7_w34_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3(0);
   bh7_w35_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3(1);
   bh7_w36_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid685: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid685_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid685_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid687_In0_c2 <= "" & bh7_w35_1_c2 & bh7_w35_2_c2 & bh7_w35_3_c2;
   bh7_w35_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3(0);
   bh7_w36_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid687: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid687_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid689_In0_c2 <= "" & bh7_w36_0_c2 & bh7_w36_1_c2 & bh7_w36_2_c2 & bh7_w36_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid689_In1_c2 <= "" & bh7_w37_0_c2;
   bh7_w36_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3(0);
   bh7_w37_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3(1);
   bh7_w38_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid689: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid689_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid689_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid691_In0_c2 <= "" & bh7_w37_1_c2 & bh7_w37_2_c2 & bh7_w37_3_c2;
   bh7_w37_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3(0);
   bh7_w38_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid691: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid691_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid693_In0_c2 <= "" & bh7_w38_0_c2 & bh7_w38_1_c2 & bh7_w38_2_c2 & bh7_w38_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid693_In1_c2 <= "" & bh7_w39_0_c2;
   bh7_w38_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3(0);
   bh7_w39_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3(1);
   bh7_w40_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid693: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid693_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid693_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid695_In0_c2 <= "" & bh7_w39_1_c2 & bh7_w39_2_c2 & bh7_w39_3_c2;
   bh7_w39_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3(0);
   bh7_w40_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid695: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid695_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid697_In0_c2 <= "" & bh7_w40_0_c2 & bh7_w40_1_c2 & bh7_w40_2_c2 & bh7_w40_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid697_In1_c2 <= "" & bh7_w41_0_c2;
   bh7_w40_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3(0);
   bh7_w41_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3(1);
   bh7_w42_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid697: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid697_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid697_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid699_In0_c2 <= "" & bh7_w41_1_c2 & bh7_w41_2_c2 & bh7_w41_3_c2;
   bh7_w41_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3(0);
   bh7_w42_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid699: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid699_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid701_In0_c2 <= "" & bh7_w42_0_c2 & bh7_w42_1_c2 & bh7_w42_2_c2 & bh7_w42_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid701_In1_c2 <= "" & bh7_w43_0_c2;
   bh7_w42_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3(0);
   bh7_w43_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3(1);
   bh7_w44_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid701: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid701_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid701_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid703_In0_c2 <= "" & bh7_w43_1_c2 & bh7_w43_2_c2 & bh7_w43_3_c2;
   bh7_w43_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3(0);
   bh7_w44_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid703: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid703_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid705_In0_c2 <= "" & bh7_w44_0_c2 & bh7_w44_1_c2 & bh7_w44_2_c2 & bh7_w44_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid705_In1_c2 <= "" & bh7_w45_0_c2;
   bh7_w44_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3(0);
   bh7_w45_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3(1);
   bh7_w46_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid705: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid705_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid705_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid707_In0_c2 <= "" & bh7_w45_1_c2 & bh7_w45_2_c2 & bh7_w45_3_c2;
   bh7_w45_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3(0);
   bh7_w46_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid707: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid707_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid709_In0_c2 <= "" & bh7_w46_0_c2 & bh7_w46_1_c2 & bh7_w46_2_c2 & bh7_w46_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid709_In1_c2 <= "" & bh7_w47_0_c2;
   bh7_w46_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3(0);
   bh7_w47_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3(1);
   bh7_w48_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid709: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid709_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid709_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid711_In0_c2 <= "" & bh7_w47_1_c2 & bh7_w47_2_c2 & bh7_w47_3_c2;
   bh7_w47_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3(0);
   bh7_w48_6_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid711: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid711_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid713_In0_c2 <= "" & bh7_w48_4_c2 & bh7_w48_0_c2 & bh7_w48_1_c2 & bh7_w48_2_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c1 <= "" & bh7_w49_5_c1;
   bh7_w48_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3(0);
   bh7_w49_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3(1);
   bh7_w50_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid713: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid713_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid715_In0_c2 <= "" & bh7_w49_0_c2 & bh7_w49_1_c2 & bh7_w49_2_c2 & bh7_w49_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c1 <= "" & bh7_w50_6_c1;
   bh7_w49_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3(0);
   bh7_w50_8_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3(1);
   bh7_w51_11_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid715: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid715_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid717_In0_c2 <= "" & bh7_w50_0_c2 & bh7_w50_1_c2 & bh7_w50_2_c2 & bh7_w50_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c1 <= "" & bh7_w51_10_c1;
   bh7_w50_9_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3(0);
   bh7_w51_12_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3(1);
   bh7_w52_12_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid717: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid717_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid719_In0_c2 <= "" & bh7_w51_0_c2 & bh7_w51_1_c2 & bh7_w51_3_c2 & bh7_w51_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c1 <= "" & bh7_w52_11_c1;
   bh7_w51_13_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3(0);
   bh7_w52_13_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3(1);
   bh7_w53_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid719: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid719_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid721_In0_c2 <= "" & bh7_w52_0_c2 & bh7_w52_1_c2 & bh7_w52_3_c2 & bh7_w52_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid721_In1_c2 <= "" & bh7_w53_14_c2;
   bh7_w52_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3(0);
   bh7_w53_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3(1);
   bh7_w54_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid721: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid721_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid721_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid723_In0_c2 <= "" & bh7_w53_0_c2 & bh7_w53_1_c2 & bh7_w53_3_c2 & bh7_w53_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid723_In1_c2 <= "" & bh7_w54_15_c2;
   bh7_w53_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3(0);
   bh7_w54_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3(1);
   bh7_w55_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid723: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid723_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid723_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid725_In0_c2 <= "" & bh7_w54_0_c2 & bh7_w54_1_c2 & bh7_w54_4_c2 & bh7_w54_5_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid725_In1_c2 <= "" & bh7_w55_17_c2;
   bh7_w54_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3(0);
   bh7_w55_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3(1);
   bh7_w56_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid725: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid725_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid725_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid727_In0_c2 <= "" & bh7_w55_0_c2 & bh7_w55_1_c2 & bh7_w55_4_c2 & bh7_w55_5_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid727_In1_c2 <= "" & bh7_w56_15_c2;
   bh7_w55_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3(0);
   bh7_w56_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3(1);
   bh7_w57_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid727: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid727_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid727_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c2 <= "" & bh7_w56_0_c2 & bh7_w56_1_c2 & bh7_w56_3_c2 & bh7_w56_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid729_In1_c3 <= "" & bh7_w57_20_c3;
   bh7_w56_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3(0);
   bh7_w57_22_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3(1);
   bh7_w58_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid729: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid729_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_copy730_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_copy730_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c2 <= "" & bh7_w57_0_c2 & bh7_w57_1_c2 & bh7_w57_4_c2 & bh7_w57_5_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid731_In1_c3 <= "" & bh7_w58_19_c3;
   bh7_w57_23_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3(0);
   bh7_w58_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3(1);
   bh7_w59_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid731: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid731_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_copy732_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_copy732_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid733_In0_c2 <= "" & bh7_w58_0_c2 & bh7_w58_3_c2 & bh7_w58_4_c2;
   bh7_w58_22_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3(0);
   bh7_w59_19_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid733: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid733_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c3; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid735_In0_c3 <= "" & bh7_w59_16_c3 & bh7_w59_17_c3 & bh7_w59_0_c3 & bh7_w59_2_c3 & bh7_w59_3_c3 & bh7_w59_4_c3;
   bh7_w59_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3(0);
   bh7_w60_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3(1);
   bh7_w61_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3(2);
   Compressor_6_3_Freq800_uid334_uid735: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid735_In0_c3,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_copy736_c3);
   Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_copy736_c3; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid737_In0_c3 <= "" & bh7_w60_19_c3 & bh7_w60_0_c3 & bh7_w60_3_c3 & bh7_w60_4_c3 & bh7_w60_5_c3;
   bh7_w60_21_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3(0);
   bh7_w61_21_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3(1);
   bh7_w62_17_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3(2);
   Compressor_5_3_Freq800_uid400_uid737: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid737_In0_c3,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_copy738_c3);
   Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_copy738_c3; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid739_In0_c3 <= "" & bh7_w61_18_c3 & bh7_w61_19_c3 & bh7_w61_0_c3 & bh7_w61_3_c3 & bh7_w61_4_c3 & bh7_w61_5_c3;
   bh7_w61_22_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3(0);
   bh7_w62_18_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3(1);
   bh7_w63_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3(2);
   Compressor_6_3_Freq800_uid334_uid739: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid739_In0_c3,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_copy740_c3);
   Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_copy740_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid741_In0_c3 <= "" & bh7_w62_16_c3 & bh7_w62_0_c3 & bh7_w62_2_c3 & bh7_w62_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid741_In1_c3 <= "" & bh7_w63_19_c3;
   bh7_w62_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3(0);
   bh7_w63_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3(1);
   bh7_w64_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid741: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid741_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid741_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_copy742_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_copy742_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid743_In0_c2 <= "" & bh7_w63_0_c2 & bh7_w63_3_c2 & bh7_w63_4_c2;
   bh7_w63_22_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3(0);
   bh7_w64_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid743: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid743_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c3; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid745_In0_c3 <= "" & bh7_w64_18_c3 & bh7_w64_19_c3 & bh7_w64_0_c3 & bh7_w64_3_c3 & bh7_w64_4_c3 & bh7_w64_5_c3;
   bh7_w64_22_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3(0);
   bh7_w65_16_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3(1);
   bh7_w66_19_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3(2);
   Compressor_6_3_Freq800_uid334_uid745: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid745_In0_c3,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_copy746_c3);
   Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_copy746_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid747_In0_c3 <= "" & bh7_w65_15_c3 & bh7_w65_0_c3 & bh7_w65_2_c3 & bh7_w65_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid747_In1_c3 <= "" & bh7_w66_18_c3;
   bh7_w65_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3(0);
   bh7_w66_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3(1);
   bh7_w67_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid747: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid747_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid747_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_copy748_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_copy748_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid749_In0_c2 <= "" & bh7_w66_0_c2 & bh7_w66_3_c2 & bh7_w66_4_c2;
   bh7_w66_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3(0);
   bh7_w67_18_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid749: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid749_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid751_In0_c3 <= "" & bh7_w67_15_c3 & bh7_w67_16_c3 & bh7_w67_0_c3 & bh7_w67_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid751_In1_c3 <= "" & bh7_w68_19_c3;
   bh7_w67_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3(0);
   bh7_w68_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3(1);
   bh7_w69_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid751: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid751_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid751_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_copy752_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_copy752_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid753_In0_c2 <= "" & bh7_w68_0_c2 & bh7_w68_2_c2 & bh7_w68_3_c2;
   bh7_w68_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3(0);
   bh7_w69_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid753: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid753_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid755_In0_c3 <= "" & bh7_w69_15_c3 & bh7_w69_0_c3 & bh7_w69_3_c3 & bh7_w69_4_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid755_In1_c3 <= "" & bh7_w70_18_c3;
   bh7_w69_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3(0);
   bh7_w70_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3(1);
   bh7_w71_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid755: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid755_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid755_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_copy756_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_copy756_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid757_In0_c3 <= "" & bh7_w70_19_c3 & bh7_w70_0_c3 & bh7_w70_3_c3 & bh7_w70_4_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid757_In1_c3 <= "" & bh7_w71_15_c3;
   bh7_w70_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3(0);
   bh7_w71_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3(1);
   bh7_w72_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid757: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid757_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid757_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_copy758_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_copy758_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid759_In0_c2 <= "" & bh7_w71_0_c2 & bh7_w71_2_c2 & bh7_w71_3_c2;
   bh7_w71_18_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3(0);
   bh7_w72_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid759: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid759_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid761_In0_c3 <= "" & bh7_w72_18_c3 & bh7_w72_19_c3 & bh7_w72_0_c3 & bh7_w72_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid761_In1_c3 <= "" & bh7_w73_15_c3;
   bh7_w72_22_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3(0);
   bh7_w73_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3(1);
   bh7_w74_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid761: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid761_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid761_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_copy762_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_copy762_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid763_In0_c2 <= "" & bh7_w73_0_c2 & bh7_w73_3_c2 & bh7_w73_4_c2;
   bh7_w73_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3(0);
   bh7_w74_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid763: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid763_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid765_In0_c3 <= "" & bh7_w74_18_c3 & bh7_w74_0_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c2 <= "" & bh7_w75_1_c2;
   bh7_w74_22_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3(0);
   bh7_w75_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3(1);
   bh7_w76_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid765: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid765_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_copy766_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_copy766_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid767_In0_c3 <= "" & bh7_w74_2_c3 & bh7_w74_3_c3 & bh7_w74_19_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid767_In1_c3 <= "" & bh7_w75_2_c3 & bh7_w75_14_c3;
   bh7_w74_23_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3(0);
   bh7_w75_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3(1);
   bh7_w76_20_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid767: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid767_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid767_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_copy768_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_copy768_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid769_In0_c3 <= "" & bh7_w76_1_c3 & bh7_w76_2_c3 & bh7_w76_18_c3 & bh7_w76_17_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c0 <= "" & "0";
   bh7_w76_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3(0);
   bh7_w77_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3(1);
   bh7_w78_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid769: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid769_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_copy770_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_copy770_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid771_In0_c3 <= "" & bh7_w77_0_c3 & bh7_w77_1_c3 & bh7_w77_14_c3;
   bh7_w77_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3(0);
   bh7_w78_20_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid771: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid771_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_copy772_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_copy772_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid773_In0_c3 <= "" & bh7_w78_0_c3 & bh7_w78_1_c3 & bh7_w78_18_c3 & bh7_w78_17_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c0 <= "" & "0";
   bh7_w78_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3(0);
   bh7_w79_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3(1);
   bh7_w80_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid773: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid773_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_copy774_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_copy774_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid775_In0_c3 <= "" & bh7_w79_0_c3 & bh7_w79_1_c3 & bh7_w79_14_c3;
   bh7_w79_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3(0);
   bh7_w80_20_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid775: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid775_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_copy776_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_copy776_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid777_In0_c3 <= "" & bh7_w80_0_c3 & bh7_w80_1_c3 & bh7_w80_18_c3 & bh7_w80_17_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c0 <= "" & "0";
   bh7_w80_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3(0);
   bh7_w81_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3(1);
   bh7_w82_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid777: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid777_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_copy778_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_copy778_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid779_In0_c3 <= "" & bh7_w81_0_c3 & bh7_w81_1_c3 & bh7_w81_14_c3;
   bh7_w81_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3(0);
   bh7_w82_20_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid779: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid779_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_copy780_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_copy780_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid781_In0_c3 <= "" & bh7_w82_18_c3 & bh7_w82_0_c3 & bh7_w82_17_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid781_In1_c3 <= "" & bh7_w83_14_c3 & bh7_w83_0_c3;
   bh7_w82_21_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3(0);
   bh7_w83_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3(1);
   bh7_w84_19_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid781: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid781_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid781_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_copy782_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_copy782_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid783_In0_c3 <= "" & bh7_w84_17_c3 & bh7_w84_18_c3 & bh7_w84_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid783_In1_c3 <= "" & bh7_w85_15_c3 & bh7_w85_0_c3;
   bh7_w84_20_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3(0);
   bh7_w85_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3(1);
   bh7_w86_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid783: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid783_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid783_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_copy784_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_copy784_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid785_In0_c3 <= "" & bh7_w86_15_c3 & bh7_w86_16_c3 & bh7_w86_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid785_In1_c3 <= "" & bh7_w87_16_c3 & bh7_w87_0_c3;
   bh7_w86_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3(0);
   bh7_w87_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3(1);
   bh7_w88_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid785: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid785_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid785_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_copy786_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_copy786_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid787_In0_c3 <= "" & bh7_w88_15_c3 & bh7_w88_16_c3 & bh7_w88_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid787_In1_c3 <= "" & bh7_w89_14_c3 & bh7_w89_0_c3;
   bh7_w88_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3(0);
   bh7_w89_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3(1);
   bh7_w90_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid787: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid787_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid787_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_copy788_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_copy788_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid789_In0_c3 <= "" & bh7_w90_15_c3 & bh7_w90_16_c3 & bh7_w90_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid789_In1_c3 <= "" & bh7_w91_15_c3 & bh7_w91_0_c3;
   bh7_w90_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3(0);
   bh7_w91_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3(1);
   bh7_w92_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid789: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid789_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid789_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_copy790_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_copy790_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid791_In0_c3 <= "" & bh7_w92_14_c3 & bh7_w92_0_c3 & "0";
   bh7_w92_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3(0);
   bh7_w93_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid791: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid791_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_copy792_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_copy792_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid793_In0_c3 <= "" & bh7_w93_15_c3 & bh7_w93_16_c3 & bh7_w93_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid793_In1_c3 <= "" & bh7_w94_15_c3 & bh7_w94_0_c3;
   bh7_w93_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3(0);
   bh7_w94_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3(1);
   bh7_w95_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid793: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid793_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid793_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_copy794_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_copy794_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid795_In0_c3 <= "" & bh7_w95_14_c3 & bh7_w95_0_c3 & "0";
   bh7_w95_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3(0);
   bh7_w96_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid795: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid795_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_copy796_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_copy796_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid797_In0_c3 <= "" & bh7_w96_15_c3 & bh7_w96_16_c3 & bh7_w96_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid797_In1_c3 <= "" & bh7_w97_15_c3 & bh7_w97_0_c3;
   bh7_w96_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3(0);
   bh7_w97_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3(1);
   bh7_w98_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid797: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid797_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid797_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_copy798_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_copy798_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid799_In0_c3 <= "" & bh7_w98_14_c3 & bh7_w98_0_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid799_In1_c3 <= "" & bh7_w99_14_c3 & bh7_w99_15_c3;
   bh7_w98_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3(0);
   bh7_w99_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3(1);
   bh7_w100_13_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid799: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid799_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid799_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_copy800_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_copy800_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid801_In0_c3 <= "" & bh7_w102_9_c3 & bh7_w102_10_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid801_In1_c3 <= "" & bh7_w103_9_c3;
   bh7_w102_11_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3(0);
   bh7_w103_10_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3(1);
   bh7_w104_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid801: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid801_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid801_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_copy802_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_copy802_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid803_In0_c3 <= "" & bh7_w105_6_c3 & bh7_w105_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c0 <= "" & "0";
   bh7_w105_8_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_c3(0);
   Compressor_14_3_Freq800_uid326_uid803: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid803_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_copy804_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_copy804_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid805_In0_c3 <= "" & bh7_w19_3_c3 & bh7_w19_2_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid805_In1_c3 <= "" & bh7_w20_2_c3;
   bh7_w19_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3(0);
   bh7_w20_3_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3(1);
   bh7_w21_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid805: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid805_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid805_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_copy806_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_copy806_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid807_In0_c3 <= "" & bh7_w21_3_c3 & bh7_w21_2_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid807_In1_c3 <= "" & bh7_w22_2_c3;
   bh7_w21_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3(0);
   bh7_w22_3_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3(1);
   bh7_w23_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid807: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid807_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid807_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_copy808_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_copy808_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid809_In0_c3 <= "" & bh7_w23_3_c3 & bh7_w23_2_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid809_In1_c3 <= "" & bh7_w24_4_c3 & bh7_w24_3_c3;
   bh7_w23_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3(0);
   bh7_w24_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3(1);
   bh7_w25_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid809: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid809_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid809_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_copy810_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_copy810_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid811_In0_c3 <= "" & bh7_w25_2_c3 & bh7_w25_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid811_In1_c3 <= "" & bh7_w26_4_c3 & bh7_w26_3_c3;
   bh7_w25_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3(0);
   bh7_w26_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3(1);
   bh7_w27_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid811: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid811_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid811_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_copy812_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_copy812_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid813_In0_c3 <= "" & bh7_w27_2_c3 & bh7_w27_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid813_In1_c3 <= "" & bh7_w28_4_c3 & bh7_w28_3_c3;
   bh7_w27_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3(0);
   bh7_w28_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3(1);
   bh7_w29_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid813: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid813_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid813_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_copy814_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_copy814_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid815_In0_c3 <= "" & bh7_w29_2_c3 & bh7_w29_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid815_In1_c3 <= "" & bh7_w30_4_c3 & bh7_w30_3_c3;
   bh7_w29_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3(0);
   bh7_w30_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3(1);
   bh7_w31_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid815: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid815_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid815_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_copy816_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_copy816_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid817_In0_c3 <= "" & bh7_w31_2_c3 & bh7_w31_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid817_In1_c3 <= "" & bh7_w32_4_c3 & bh7_w32_3_c3;
   bh7_w31_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3(0);
   bh7_w32_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3(1);
   bh7_w33_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid817: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid817_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid817_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_copy818_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_copy818_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid819_In0_c3 <= "" & bh7_w33_2_c3 & bh7_w33_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid819_In1_c3 <= "" & bh7_w34_5_c3 & bh7_w34_4_c3;
   bh7_w33_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3(0);
   bh7_w34_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3(1);
   bh7_w35_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid819: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid819_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid819_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_copy820_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_copy820_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid821_In0_c3 <= "" & bh7_w35_5_c3 & bh7_w35_4_c3 & "0";
   bh7_w35_7_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3(0);
   bh7_w36_7_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid821: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid821_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_copy822_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_copy822_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid823_In0_c3 <= "" & bh7_w36_6_c3 & bh7_w36_5_c3 & bh7_w36_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid823_In1_c3 <= "" & bh7_w37_5_c3 & bh7_w37_4_c3;
   bh7_w36_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3(0);
   bh7_w37_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3(1);
   bh7_w38_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid823: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid823_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid823_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_copy824_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_copy824_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid825_In0_c3 <= "" & bh7_w38_6_c3 & bh7_w38_5_c3 & bh7_w38_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid825_In1_c3 <= "" & bh7_w39_5_c3 & bh7_w39_4_c3;
   bh7_w38_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3(0);
   bh7_w39_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3(1);
   bh7_w40_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid825: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid825_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid825_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_copy826_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_copy826_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid827_In0_c3 <= "" & bh7_w40_6_c3 & bh7_w40_5_c3 & bh7_w40_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid827_In1_c3 <= "" & bh7_w41_5_c3 & bh7_w41_4_c3;
   bh7_w40_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3(0);
   bh7_w41_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3(1);
   bh7_w42_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid827: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid827_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid827_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_copy828_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_copy828_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid829_In0_c3 <= "" & bh7_w42_6_c3 & bh7_w42_5_c3 & bh7_w42_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid829_In1_c3 <= "" & bh7_w43_5_c3 & bh7_w43_4_c3;
   bh7_w42_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3(0);
   bh7_w43_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3(1);
   bh7_w44_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid829: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid829_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid829_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_copy830_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_copy830_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid831_In0_c3 <= "" & bh7_w44_6_c3 & bh7_w44_5_c3 & bh7_w44_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid831_In1_c3 <= "" & bh7_w45_5_c3 & bh7_w45_4_c3;
   bh7_w44_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3(0);
   bh7_w45_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3(1);
   bh7_w46_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid831: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid831_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid831_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_copy832_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_copy832_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid833_In0_c3 <= "" & bh7_w46_6_c3 & bh7_w46_5_c3 & bh7_w46_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid833_In1_c3 <= "" & bh7_w47_5_c3 & bh7_w47_4_c3;
   bh7_w46_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3(0);
   bh7_w47_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3(1);
   bh7_w48_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid833: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid833_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid833_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_copy834_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_copy834_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid835_In0_c3 <= "" & bh7_w48_3_c3 & bh7_w48_7_c3 & bh7_w48_6_c3 & bh7_w48_5_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid835_In1_c3 <= "" & bh7_w49_7_c3;
   bh7_w48_9_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3(0);
   bh7_w49_8_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3(1);
   bh7_w50_10_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid835: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid835_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid835_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_copy836_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_copy836_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid837_In0_c3 <= "" & bh7_w50_9_c3 & bh7_w50_8_c3 & bh7_w50_7_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid837_In1_c3 <= "" & bh7_w51_13_c3 & bh7_w51_12_c3;
   bh7_w50_11_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3(0);
   bh7_w51_14_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3(1);
   bh7_w52_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid837: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid837_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid837_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_copy838_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_copy838_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid839_In0_c3 <= "" & bh7_w52_14_c3 & bh7_w52_13_c3 & bh7_w52_12_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid839_In1_c3 <= "" & bh7_w53_17_c3 & bh7_w53_16_c3;
   bh7_w52_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3(0);
   bh7_w53_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3(1);
   bh7_w54_19_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid839: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid839_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid839_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_copy840_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_copy840_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid841_In0_c3 <= "" & bh7_w54_18_c3 & bh7_w54_17_c3 & bh7_w54_16_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid841_In1_c3 <= "" & bh7_w55_19_c3 & bh7_w55_20_c3;
   bh7_w54_20_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3(0);
   bh7_w55_21_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3(1);
   bh7_w56_19_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid841: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid841_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid841_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_copy842_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_copy842_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid843_In0_c3 <= "" & bh7_w56_16_c3 & bh7_w56_17_c3 & bh7_w56_18_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid843_In1_c3 <= "" & bh7_w57_21_c3 & bh7_w57_22_c3;
   bh7_w56_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4(0);
   bh7_w57_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4(1);
   bh7_w58_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid843: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid843_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid843_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid845_In0_c3 <= "" & bh7_w58_20_c3 & bh7_w58_21_c3 & bh7_w58_5_c3 & bh7_w58_22_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c0 <= "" & "0";
   bh7_w58_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4(0);
   bh7_w59_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4(1);
   bh7_w60_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid845: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid845_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid847_In0_c3 <= "" & bh7_w59_18_c3 & bh7_w59_20_c3 & bh7_w59_19_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid847_In1_c3 <= "" & bh7_w60_20_c3 & bh7_w60_21_c3;
   bh7_w59_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4(0);
   bh7_w60_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4(1);
   bh7_w61_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid847: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid847_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid847_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid849_In0_c3 <= "" & bh7_w61_20_c3 & bh7_w61_21_c3 & bh7_w61_22_c3;
   bh7_w61_24_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4(0);
   bh7_w62_20_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid849: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid849_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid851_In0_c3 <= "" & bh7_w62_17_c3 & bh7_w62_18_c3 & bh7_w62_19_c3 & bh7_w62_4_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid851_In1_c3 <= "" & bh7_w63_20_c3;
   bh7_w62_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4(0);
   bh7_w63_23_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4(1);
   bh7_w64_23_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid851: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid851_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid851_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid853_In0_c3 <= "" & bh7_w63_21_c3 & bh7_w63_5_c3 & bh7_w63_22_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c0 <= "" & "0" & "0";
   bh7_w63_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4(0);
   bh7_w64_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4(1);
   bh7_w65_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid853: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid853_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid855_In0_c3 <= "" & bh7_w64_20_c3 & bh7_w64_22_c3 & bh7_w64_21_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid855_In1_c3 <= "" & bh7_w65_16_c3 & bh7_w65_17_c3;
   bh7_w64_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4(0);
   bh7_w65_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4(1);
   bh7_w66_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid855: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid855_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid855_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid857_In0_c3 <= "" & bh7_w66_19_c3 & bh7_w66_20_c3 & bh7_w66_21_c3;
   bh7_w66_23_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4(0);
   bh7_w67_20_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid857: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid857_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid859_In0_c3 <= "" & bh7_w67_17_c3 & bh7_w67_19_c3 & bh7_w67_4_c3 & bh7_w67_18_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid859_In1_c3 <= "" & bh7_w68_20_c3;
   bh7_w67_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4(0);
   bh7_w68_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4(1);
   bh7_w69_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid859: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid859_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid859_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid861_In0_c3 <= "" & bh7_w69_16_c3 & bh7_w69_18_c3 & bh7_w69_17_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid861_In1_c3 <= "" & bh7_w70_20_c3 & bh7_w70_21_c3;
   bh7_w69_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4(0);
   bh7_w70_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4(1);
   bh7_w71_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid861: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid861_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid861_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid863_In0_c3 <= "" & bh7_w71_16_c3 & bh7_w71_17_c3 & bh7_w71_18_c3;
   bh7_w71_20_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4(0);
   bh7_w72_23_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid863: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid863_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid865_In0_c3 <= "" & bh7_w72_20_c3 & bh7_w72_22_c3 & bh7_w72_4_c3 & bh7_w72_21_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid865_In1_c3 <= "" & bh7_w73_16_c3;
   bh7_w72_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4(0);
   bh7_w73_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4(1);
   bh7_w74_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid865: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid865_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid865_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid867_In0_c3 <= "" & bh7_w74_20_c3 & bh7_w74_22_c3 & bh7_w74_21_c3 & bh7_w74_23_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid867_In1_c3 <= "" & bh7_w75_15_c3;
   bh7_w74_25_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4(0);
   bh7_w75_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4(1);
   bh7_w76_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid867: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid867_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid867_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid869_In0_c3 <= "" & bh7_w76_19_c3 & bh7_w76_21_c3 & bh7_w76_20_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid869_In1_c3 <= "" & bh7_w77_15_c3 & bh7_w77_16_c3;
   bh7_w76_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4(0);
   bh7_w77_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4(1);
   bh7_w78_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid869: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid869_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid869_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid871_In0_c3 <= "" & bh7_w78_19_c3 & bh7_w78_21_c3 & bh7_w78_20_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid871_In1_c3 <= "" & bh7_w79_15_c3 & bh7_w79_16_c3;
   bh7_w78_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4(0);
   bh7_w79_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4(1);
   bh7_w80_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid871: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid871_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid871_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid873_In0_c3 <= "" & bh7_w80_19_c3 & bh7_w80_21_c3 & bh7_w80_20_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid873_In1_c3 <= "" & bh7_w81_15_c3 & bh7_w81_16_c3;
   bh7_w80_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4(0);
   bh7_w81_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4(1);
   bh7_w82_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid873: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid873_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid873_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid875_In0_c3 <= "" & bh7_w82_19_c3 & bh7_w82_21_c3 & bh7_w82_20_c3;
   bh7_w82_23_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4(0);
   bh7_w83_16_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid875: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid875_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid877_In0_c3 <= "" & bh7_w84_19_c3 & bh7_w84_20_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid877_In1_c3 <= "" & bh7_w85_16_c3;
   bh7_w84_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4(0);
   bh7_w85_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4(1);
   bh7_w86_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid877: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid877_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid877_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid879_In0_c3 <= "" & bh7_w86_17_c3 & bh7_w86_18_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid879_In1_c3 <= "" & bh7_w87_17_c3;
   bh7_w86_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4(0);
   bh7_w87_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4(1);
   bh7_w88_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid879: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid879_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid879_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid881_In0_c3 <= "" & bh7_w88_17_c3 & bh7_w88_18_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid881_In1_c3 <= "" & bh7_w89_15_c3;
   bh7_w88_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4(0);
   bh7_w89_16_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4(1);
   bh7_w90_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid881: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid881_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid881_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid883_In0_c3 <= "" & bh7_w90_17_c3 & bh7_w90_18_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid883_In1_c3 <= "" & bh7_w91_16_c3;
   bh7_w90_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4(0);
   bh7_w91_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4(1);
   bh7_w92_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid883: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid883_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid883_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid885_In0_c3 <= "" & bh7_w92_15_c3 & bh7_w92_16_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid885_In1_c3 <= "" & bh7_w93_17_c3 & bh7_w93_18_c3;
   bh7_w92_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4(0);
   bh7_w93_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4(1);
   bh7_w94_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid885: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid885_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid885_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid887_In0_c3 <= "" & bh7_w95_15_c3 & bh7_w95_16_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid887_In1_c3 <= "" & bh7_w96_17_c3 & bh7_w96_18_c3;
   bh7_w95_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4(0);
   bh7_w96_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4(1);
   bh7_w97_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid887: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid887_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid887_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid889_In0_c3 <= "" & bh7_w98_15_c3 & bh7_w98_16_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid889_In1_c3 <= "" & bh7_w99_16_c3;
   bh7_w98_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4(0);
   bh7_w99_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4(1);
   bh7_w100_14_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid889: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid889_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid889_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid891_In0_c3 <= "" & bh7_w100_12_c3 & bh7_w100_13_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid891_In1_c3 <= "" & bh7_w101_11_c3;
   bh7_w100_15_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4(0);
   bh7_w101_12_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4(1);
   bh7_w102_12_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid891: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid891_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid891_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid893_In0_c3 <= "" & bh7_w104_5_c3 & bh7_w104_6_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid893_In1_c3 <= "" & bh7_w105_8_c3;
   bh7_w104_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4(0);
   bh7_w105_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4(1);
   Compressor_14_3_Freq800_uid326_uid893: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid893_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid893_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid895_In0_c3 <= "" & bh7_w21_5_c3 & bh7_w21_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid895_In1_c3 <= "" & bh7_w22_3_c3;
   bh7_w21_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4(0);
   bh7_w22_4_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4(1);
   bh7_w23_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid895: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid895_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid895_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid897_In0_c3 <= "" & bh7_w23_5_c3 & bh7_w23_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid897_In1_c3 <= "" & bh7_w24_5_c3;
   bh7_w23_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4(0);
   bh7_w24_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4(1);
   bh7_w25_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid897: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid897_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid897_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid899_In0_c3 <= "" & bh7_w25_5_c3 & bh7_w25_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid899_In1_c3 <= "" & bh7_w26_5_c3;
   bh7_w25_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4(0);
   bh7_w26_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4(1);
   bh7_w27_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid899: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid899_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid899_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid901_In0_c3 <= "" & bh7_w27_5_c3 & bh7_w27_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid901_In1_c3 <= "" & bh7_w28_5_c3;
   bh7_w27_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4(0);
   bh7_w28_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4(1);
   bh7_w29_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid901: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid901_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid901_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid903_In0_c3 <= "" & bh7_w29_5_c3 & bh7_w29_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid903_In1_c3 <= "" & bh7_w30_5_c3;
   bh7_w29_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4(0);
   bh7_w30_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4(1);
   bh7_w31_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid903: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid903_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid903_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid905_In0_c3 <= "" & bh7_w31_5_c3 & bh7_w31_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid905_In1_c3 <= "" & bh7_w32_5_c3;
   bh7_w31_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4(0);
   bh7_w32_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4(1);
   bh7_w33_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid905: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid905_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid905_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid907_In0_c3 <= "" & bh7_w33_5_c3 & bh7_w33_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid907_In1_c3 <= "" & bh7_w34_6_c3;
   bh7_w33_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4(0);
   bh7_w34_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4(1);
   bh7_w35_8_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid907: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid907_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid907_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid909_In0_c3 <= "" & bh7_w35_7_c3 & bh7_w35_6_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid909_In1_c3 <= "" & bh7_w36_8_c3 & bh7_w36_7_c3;
   bh7_w35_9_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4(0);
   bh7_w36_9_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4(1);
   bh7_w37_7_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid909: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid909_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid909_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid911_In0_c3 <= "" & bh7_w38_8_c3 & bh7_w38_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid911_In1_c3 <= "" & bh7_w39_6_c3;
   bh7_w38_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4(0);
   bh7_w39_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4(1);
   bh7_w40_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid911: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid911_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid911_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid913_In0_c3 <= "" & bh7_w40_8_c3 & bh7_w40_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid913_In1_c3 <= "" & bh7_w41_6_c3;
   bh7_w40_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4(0);
   bh7_w41_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4(1);
   bh7_w42_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid913: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid913_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid913_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid915_In0_c3 <= "" & bh7_w42_8_c3 & bh7_w42_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid915_In1_c3 <= "" & bh7_w43_6_c3;
   bh7_w42_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4(0);
   bh7_w43_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4(1);
   bh7_w44_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid915: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid915_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid915_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid917_In0_c3 <= "" & bh7_w44_8_c3 & bh7_w44_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid917_In1_c3 <= "" & bh7_w45_6_c3;
   bh7_w44_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4(0);
   bh7_w45_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4(1);
   bh7_w46_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid917: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid917_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid917_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid919_In0_c3 <= "" & bh7_w46_8_c3 & bh7_w46_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid919_In1_c3 <= "" & bh7_w47_6_c3;
   bh7_w46_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4(0);
   bh7_w47_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4(1);
   bh7_w48_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid919: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid919_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid919_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid921_In0_c3 <= "" & bh7_w48_9_c3 & bh7_w48_8_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid921_In1_c3 <= "" & bh7_w49_6_c3 & bh7_w49_8_c3;
   bh7_w48_11_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4(0);
   bh7_w49_9_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4(1);
   bh7_w50_12_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid921: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid921_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid921_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid923_In0_c3 <= "" & bh7_w50_11_c3 & bh7_w50_10_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid923_In1_c3 <= "" & bh7_w51_11_c3 & bh7_w51_14_c3;
   bh7_w50_13_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4(0);
   bh7_w51_15_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4(1);
   bh7_w52_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid923: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid923_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid923_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid925_In0_c3 <= "" & bh7_w52_16_c3 & bh7_w52_15_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid925_In1_c3 <= "" & bh7_w53_15_c3 & bh7_w53_18_c3;
   bh7_w52_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4(0);
   bh7_w53_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4(1);
   bh7_w54_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid925: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid925_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid925_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid927_In0_c3 <= "" & bh7_w54_20_c3 & bh7_w54_19_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid927_In1_c3 <= "" & bh7_w55_21_c3 & bh7_w55_18_c3;
   bh7_w54_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4(0);
   bh7_w55_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4(1);
   bh7_w56_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid927: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid927_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid927_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid929_In0_c4 <= "" & bh7_w56_19_c4 & bh7_w56_20_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid929_In1_c4 <= "" & bh7_w57_23_c4 & bh7_w57_24_c4;
   bh7_w56_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4(0);
   bh7_w57_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4(1);
   bh7_w58_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid929: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid929_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid929_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_copy930_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_copy930_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid931_In0_c4 <= "" & bh7_w58_23_c4 & bh7_w58_24_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid931_In1_c4 <= "" & bh7_w59_21_c4 & bh7_w59_22_c4;
   bh7_w58_26_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4(0);
   bh7_w59_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4(1);
   bh7_w60_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid931: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid931_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid931_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_copy932_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_copy932_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid933_In0_c4 <= "" & bh7_w60_22_c4 & bh7_w60_23_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid933_In1_c4 <= "" & bh7_w61_23_c4 & bh7_w61_24_c4;
   bh7_w60_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4(0);
   bh7_w61_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4(1);
   bh7_w62_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid933: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid933_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid933_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_copy934_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_copy934_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid935_In0_c4 <= "" & bh7_w62_20_c4 & bh7_w62_21_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid935_In1_c4 <= "" & bh7_w63_23_c4 & bh7_w63_24_c4;
   bh7_w62_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4(0);
   bh7_w63_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4(1);
   bh7_w64_26_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid935: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid935_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid935_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_copy936_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_copy936_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid937_In0_c4 <= "" & bh7_w64_23_c4 & bh7_w64_24_c4 & bh7_w64_25_c4;
   Compressor_23_3_Freq800_uid322_bh7_uid937_In1_c4 <= "" & bh7_w65_18_c4 & bh7_w65_19_c4;
   bh7_w64_27_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4(0);
   bh7_w65_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4(1);
   bh7_w66_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid937: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid937_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid937_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_copy938_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_copy938_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid939_In0_c4 <= "" & bh7_w66_22_c4 & bh7_w66_23_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid939_In1_c4 <= "" & bh7_w67_20_c4 & bh7_w67_21_c4;
   bh7_w66_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4(0);
   bh7_w67_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4(1);
   bh7_w68_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid939: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid939_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid939_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_copy940_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_copy940_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid941_In0_c4 <= "" & bh7_w68_22_c4 & bh7_w68_21_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid941_In1_c4 <= "" & bh7_w69_19_c4 & bh7_w69_20_c4;
   bh7_w68_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4(0);
   bh7_w69_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4(1);
   bh7_w70_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid941: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid941_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid941_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_copy942_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_copy942_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid943_In0_c4 <= "" & bh7_w71_19_c4 & bh7_w71_20_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid943_In1_c4 <= "" & bh7_w72_23_c4 & bh7_w72_24_c4;
   bh7_w71_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4(0);
   bh7_w72_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4(1);
   bh7_w73_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid943: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid943_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid943_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_copy944_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_copy944_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid945_In0_c4 <= "" & bh7_w73_18_c4 & bh7_w73_17_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid945_In1_c4 <= "" & bh7_w74_24_c4 & bh7_w74_25_c4;
   bh7_w73_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4(0);
   bh7_w74_26_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4(1);
   bh7_w75_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid945: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid945_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid945_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_copy946_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_copy946_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid947_In0_c4 <= "" & bh7_w75_17_c4 & bh7_w75_16_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid947_In1_c4 <= "" & bh7_w76_22_c4 & bh7_w76_23_c4;
   bh7_w75_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4(0);
   bh7_w76_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4(1);
   bh7_w77_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid947: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid947_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid947_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_copy948_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_copy948_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid949_In0_c4 <= "" & bh7_w78_22_c4 & bh7_w78_23_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid949_In1_c4 <= "" & bh7_w79_17_c4;
   bh7_w78_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4(0);
   bh7_w79_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4(1);
   bh7_w80_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid949: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid949_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid949_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_copy950_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_copy950_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid951_In0_c4 <= "" & bh7_w80_22_c4 & bh7_w80_23_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid951_In1_c4 <= "" & bh7_w81_17_c4;
   bh7_w80_25_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4(0);
   bh7_w81_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4(1);
   bh7_w82_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid951: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid951_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid951_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_copy952_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_copy952_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid953_In0_c4 <= "" & bh7_w82_22_c4 & bh7_w82_23_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid953_In1_c4 <= "" & bh7_w83_15_c4 & bh7_w83_16_c4;
   bh7_w82_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4(0);
   bh7_w83_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4(1);
   bh7_w84_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid953: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid953_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid953_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_copy954_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_copy954_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid955_In0_c4 <= "" & bh7_w86_19_c4 & bh7_w86_20_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid955_In1_c4 <= "" & bh7_w87_18_c4;
   bh7_w86_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4(0);
   bh7_w87_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4(1);
   bh7_w88_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid955: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid955_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid955_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_copy956_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_copy956_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid957_In0_c4 <= "" & bh7_w88_19_c4 & bh7_w88_20_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid957_In1_c4 <= "" & bh7_w89_16_c4;
   bh7_w88_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4(0);
   bh7_w89_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4(1);
   bh7_w90_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid957: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid957_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid957_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_copy958_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_copy958_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid959_In0_c4 <= "" & bh7_w90_19_c4 & bh7_w90_20_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid959_In1_c4 <= "" & bh7_w91_17_c4;
   bh7_w90_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4(0);
   bh7_w91_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4(1);
   bh7_w92_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid959: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid959_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid959_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_copy960_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_copy960_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid961_In0_c4 <= "" & bh7_w92_17_c4 & bh7_w92_18_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid961_In1_c4 <= "" & bh7_w93_19_c4;
   bh7_w92_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4(0);
   bh7_w93_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4(1);
   bh7_w94_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid961: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid961_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid961_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_copy962_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_copy962_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid963_In0_c4 <= "" & bh7_w94_16_c4 & bh7_w94_17_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid963_In1_c4 <= "" & bh7_w95_17_c4;
   bh7_w94_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4(0);
   bh7_w95_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4(1);
   bh7_w96_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid963: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid963_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid963_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_copy964_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_copy964_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid965_In0_c4 <= "" & bh7_w97_16_c4 & bh7_w97_17_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid965_In1_c4 <= "" & bh7_w98_17_c4;
   bh7_w97_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4(0);
   bh7_w98_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4(1);
   bh7_w99_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid965: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid965_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid965_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_copy966_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_copy966_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid967_In0_c4 <= "" & bh7_w100_14_c4 & bh7_w100_15_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid967_In1_c4 <= "" & bh7_w101_12_c4;
   bh7_w100_16_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4(0);
   bh7_w101_13_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4(1);
   bh7_w102_13_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid967: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid967_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid967_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_copy968_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_copy968_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid969_In0_c4 <= "" & bh7_w102_11_c4 & bh7_w102_12_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c3 <= "" & bh7_w103_10_c3;
   bh7_w102_14_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4(0);
   bh7_w103_11_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4(1);
   bh7_w104_8_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid969: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid969_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_copy970_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_copy970_c4; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_22_c4 <= bh7_w22_4_c4 & bh7_w21_6_c4 & bh7_w20_3_c4 & bh7_w19_4_c4 & bh7_w18_2_c4 & bh7_w17_2_c4 & bh7_w16_0_c4 & bh7_w15_0_c4 & bh7_w14_0_c4 & bh7_w13_0_c4 & bh7_w12_0_c4 & bh7_w11_0_c4 & bh7_w10_0_c4 & bh7_w9_0_c4 & bh7_w8_0_c4 & bh7_w7_0_c4 & bh7_w6_0_c4 & bh7_w5_0_c4 & bh7_w4_0_c4 & bh7_w3_0_c4 & bh7_w2_0_c4 & bh7_w1_0_c4 & bh7_w0_0_c4;

   bitheapFinalAdd_bh7_In0_c4 <= "0" & bh7_w105_9_c4 & bh7_w104_7_c4 & bh7_w103_11_c4 & bh7_w102_13_c4 & bh7_w101_13_c4 & bh7_w100_16_c4 & bh7_w99_17_c4 & bh7_w98_18_c4 & bh7_w97_18_c4 & bh7_w96_19_c4 & bh7_w95_18_c4 & bh7_w94_18_c4 & bh7_w93_20_c4 & bh7_w92_19_c4 & bh7_w91_18_c4 & bh7_w90_21_c4 & bh7_w89_17_c4 & bh7_w88_21_c4 & bh7_w87_19_c4 & bh7_w86_21_c4 & bh7_w85_17_c4 & bh7_w84_21_c4 & bh7_w83_17_c4 & bh7_w82_24_c4 & bh7_w81_18_c4 & bh7_w80_24_c4 & bh7_w79_18_c4 & bh7_w78_24_c4 & bh7_w77_17_c4 & bh7_w76_24_c4 & bh7_w75_18_c4 & bh7_w74_26_c4 & bh7_w73_19_c4 & bh7_w72_25_c4 & bh7_w71_21_c4 & bh7_w70_22_c4 & bh7_w69_21_c4 & bh7_w68_23_c4 & bh7_w67_22_c4 & bh7_w66_24_c4 & bh7_w65_20_c4 & bh7_w64_26_c4 & bh7_w63_25_c4 & bh7_w62_22_c4 & bh7_w61_25_c4 & bh7_w60_24_c4 & bh7_w59_23_c4 & bh7_w58_25_c4 & bh7_w57_25_c4 & bh7_w56_21_c4 & bh7_w55_22_c4 & bh7_w54_22_c4 & bh7_w53_19_c4 & bh7_w52_18_c4 & bh7_w51_15_c4 & bh7_w50_13_c4 & bh7_w49_9_c4 & bh7_w48_11_c4 & bh7_w47_7_c4 & bh7_w46_10_c4 & bh7_w45_7_c4 & bh7_w44_10_c4 & bh7_w43_7_c4 & bh7_w42_10_c4 & bh7_w41_7_c4 & bh7_w40_10_c4 & bh7_w39_7_c4 & bh7_w38_9_c4 & bh7_w37_6_c4 & bh7_w36_9_c4 & bh7_w35_9_c4 & bh7_w34_7_c4 & bh7_w33_7_c4 & bh7_w32_6_c4 & bh7_w31_7_c4 & bh7_w30_6_c4 & bh7_w29_7_c4 & bh7_w28_6_c4 & bh7_w27_7_c4 & bh7_w26_6_c4 & bh7_w25_7_c4 & bh7_w24_6_c4 & bh7_w23_7_c4;
   bitheapFinalAdd_bh7_In1_c4 <= "0" & "0" & bh7_w104_8_c4 & "0" & bh7_w102_14_c4 & "0" & "0" & bh7_w99_18_c4 & "0" & "0" & bh7_w96_20_c4 & "0" & bh7_w94_19_c4 & "0" & bh7_w92_20_c4 & "0" & bh7_w90_22_c4 & "0" & bh7_w88_22_c4 & "0" & "0" & "0" & bh7_w84_22_c4 & "0" & bh7_w82_25_c4 & "0" & bh7_w80_25_c4 & "0" & "0" & bh7_w77_18_c4 & "0" & bh7_w75_19_c4 & "0" & bh7_w73_20_c4 & "0" & "0" & bh7_w70_23_c4 & "0" & bh7_w68_24_c4 & "0" & bh7_w66_25_c4 & "0" & bh7_w64_27_c4 & "0" & bh7_w62_23_c4 & "0" & bh7_w60_25_c4 & "0" & bh7_w58_26_c4 & "0" & bh7_w56_22_c4 & "0" & bh7_w54_21_c4 & "0" & bh7_w52_17_c4 & "0" & bh7_w50_12_c4 & "0" & bh7_w48_10_c4 & "0" & bh7_w46_9_c4 & "0" & bh7_w44_9_c4 & "0" & bh7_w42_9_c4 & "0" & bh7_w40_9_c4 & "0" & "0" & bh7_w37_7_c4 & "0" & bh7_w35_8_c4 & "0" & bh7_w33_6_c4 & "0" & bh7_w31_6_c4 & "0" & bh7_w29_6_c4 & "0" & bh7_w27_6_c4 & "0" & bh7_w25_6_c4 & "0" & bh7_w23_6_c4;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_84_Freq800_uid972
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c4,
                 Y => bitheapFinalAdd_bh7_In1_c4,
                 R => bitheapFinalAdd_bh7_Out_c33);
   bitheapResult_bh7_c33 <= bitheapFinalAdd_bh7_Out_c33(82 downto 0) & tmp_bitheapResult_bh7_22_c33;
   R <= bitheapResult_bh7_c33(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_65_Freq800_uid975
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq800_uid975 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq800_uid975 is
signal Cin_1_c34, Cin_1_c35 :  std_logic;
signal X_1_c33, X_1_c34, X_1_c35 :  std_logic_vector(3 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9, Y_1_c10, Y_1_c11, Y_1_c12, Y_1_c13, Y_1_c14, Y_1_c15, Y_1_c16, Y_1_c17, Y_1_c18, Y_1_c19, Y_1_c20, Y_1_c21, Y_1_c22, Y_1_c23, Y_1_c24, Y_1_c25, Y_1_c26, Y_1_c27, Y_1_c28, Y_1_c29, Y_1_c30, Y_1_c31, Y_1_c32, Y_1_c33, Y_1_c34, Y_1_c35 :  std_logic_vector(3 downto 0);
signal S_1_c35 :  std_logic_vector(3 downto 0);
signal R_1_c35, R_1_c36, R_1_c37, R_1_c38, R_1_c39, R_1_c40, R_1_c41, R_1_c42, R_1_c43, R_1_c44, R_1_c45, R_1_c46, R_1_c47, R_1_c48, R_1_c49, R_1_c50, R_1_c51, R_1_c52, R_1_c53, R_1_c54, R_1_c55, R_1_c56 :  std_logic_vector(2 downto 0);
signal Cin_2_c35, Cin_2_c36 :  std_logic;
signal X_2_c33, X_2_c34, X_2_c35, X_2_c36 :  std_logic_vector(3 downto 0);
signal Y_2_c0, Y_2_c1, Y_2_c2, Y_2_c3, Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7, Y_2_c8, Y_2_c9, Y_2_c10, Y_2_c11, Y_2_c12, Y_2_c13, Y_2_c14, Y_2_c15, Y_2_c16, Y_2_c17, Y_2_c18, Y_2_c19, Y_2_c20, Y_2_c21, Y_2_c22, Y_2_c23, Y_2_c24, Y_2_c25, Y_2_c26, Y_2_c27, Y_2_c28, Y_2_c29, Y_2_c30, Y_2_c31, Y_2_c32, Y_2_c33, Y_2_c34, Y_2_c35, Y_2_c36 :  std_logic_vector(3 downto 0);
signal S_2_c36 :  std_logic_vector(3 downto 0);
signal R_2_c36, R_2_c37, R_2_c38, R_2_c39, R_2_c40, R_2_c41, R_2_c42, R_2_c43, R_2_c44, R_2_c45, R_2_c46, R_2_c47, R_2_c48, R_2_c49, R_2_c50, R_2_c51, R_2_c52, R_2_c53, R_2_c54, R_2_c55, R_2_c56 :  std_logic_vector(2 downto 0);
signal Cin_3_c36, Cin_3_c37 :  std_logic;
signal X_3_c33, X_3_c34, X_3_c35, X_3_c36, X_3_c37 :  std_logic_vector(3 downto 0);
signal Y_3_c0, Y_3_c1, Y_3_c2, Y_3_c3, Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8, Y_3_c9, Y_3_c10, Y_3_c11, Y_3_c12, Y_3_c13, Y_3_c14, Y_3_c15, Y_3_c16, Y_3_c17, Y_3_c18, Y_3_c19, Y_3_c20, Y_3_c21, Y_3_c22, Y_3_c23, Y_3_c24, Y_3_c25, Y_3_c26, Y_3_c27, Y_3_c28, Y_3_c29, Y_3_c30, Y_3_c31, Y_3_c32, Y_3_c33, Y_3_c34, Y_3_c35, Y_3_c36, Y_3_c37 :  std_logic_vector(3 downto 0);
signal S_3_c37 :  std_logic_vector(3 downto 0);
signal R_3_c37, R_3_c38, R_3_c39, R_3_c40, R_3_c41, R_3_c42, R_3_c43, R_3_c44, R_3_c45, R_3_c46, R_3_c47, R_3_c48, R_3_c49, R_3_c50, R_3_c51, R_3_c52, R_3_c53, R_3_c54, R_3_c55, R_3_c56 :  std_logic_vector(2 downto 0);
signal Cin_4_c37, Cin_4_c38 :  std_logic;
signal X_4_c33, X_4_c34, X_4_c35, X_4_c36, X_4_c37, X_4_c38 :  std_logic_vector(3 downto 0);
signal Y_4_c0, Y_4_c1, Y_4_c2, Y_4_c3, Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9, Y_4_c10, Y_4_c11, Y_4_c12, Y_4_c13, Y_4_c14, Y_4_c15, Y_4_c16, Y_4_c17, Y_4_c18, Y_4_c19, Y_4_c20, Y_4_c21, Y_4_c22, Y_4_c23, Y_4_c24, Y_4_c25, Y_4_c26, Y_4_c27, Y_4_c28, Y_4_c29, Y_4_c30, Y_4_c31, Y_4_c32, Y_4_c33, Y_4_c34, Y_4_c35, Y_4_c36, Y_4_c37, Y_4_c38 :  std_logic_vector(3 downto 0);
signal S_4_c38 :  std_logic_vector(3 downto 0);
signal R_4_c38, R_4_c39, R_4_c40, R_4_c41, R_4_c42, R_4_c43, R_4_c44, R_4_c45, R_4_c46, R_4_c47, R_4_c48, R_4_c49, R_4_c50, R_4_c51, R_4_c52, R_4_c53, R_4_c54, R_4_c55, R_4_c56 :  std_logic_vector(2 downto 0);
signal Cin_5_c38, Cin_5_c39 :  std_logic;
signal X_5_c33, X_5_c34, X_5_c35, X_5_c36, X_5_c37, X_5_c38, X_5_c39 :  std_logic_vector(3 downto 0);
signal Y_5_c0, Y_5_c1, Y_5_c2, Y_5_c3, Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13, Y_5_c14, Y_5_c15, Y_5_c16, Y_5_c17, Y_5_c18, Y_5_c19, Y_5_c20, Y_5_c21, Y_5_c22, Y_5_c23, Y_5_c24, Y_5_c25, Y_5_c26, Y_5_c27, Y_5_c28, Y_5_c29, Y_5_c30, Y_5_c31, Y_5_c32, Y_5_c33, Y_5_c34, Y_5_c35, Y_5_c36, Y_5_c37, Y_5_c38, Y_5_c39 :  std_logic_vector(3 downto 0);
signal S_5_c39 :  std_logic_vector(3 downto 0);
signal R_5_c39, R_5_c40, R_5_c41, R_5_c42, R_5_c43, R_5_c44, R_5_c45, R_5_c46, R_5_c47, R_5_c48, R_5_c49, R_5_c50, R_5_c51, R_5_c52, R_5_c53, R_5_c54, R_5_c55, R_5_c56 :  std_logic_vector(2 downto 0);
signal Cin_6_c39, Cin_6_c40 :  std_logic;
signal X_6_c33, X_6_c34, X_6_c35, X_6_c36, X_6_c37, X_6_c38, X_6_c39, X_6_c40 :  std_logic_vector(3 downto 0);
signal Y_6_c0, Y_6_c1, Y_6_c2, Y_6_c3, Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11, Y_6_c12, Y_6_c13, Y_6_c14, Y_6_c15, Y_6_c16, Y_6_c17, Y_6_c18, Y_6_c19, Y_6_c20, Y_6_c21, Y_6_c22, Y_6_c23, Y_6_c24, Y_6_c25, Y_6_c26, Y_6_c27, Y_6_c28, Y_6_c29, Y_6_c30, Y_6_c31, Y_6_c32, Y_6_c33, Y_6_c34, Y_6_c35, Y_6_c36, Y_6_c37, Y_6_c38, Y_6_c39, Y_6_c40 :  std_logic_vector(3 downto 0);
signal S_6_c40 :  std_logic_vector(3 downto 0);
signal R_6_c40, R_6_c41, R_6_c42, R_6_c43, R_6_c44, R_6_c45, R_6_c46, R_6_c47, R_6_c48, R_6_c49, R_6_c50, R_6_c51, R_6_c52, R_6_c53, R_6_c54, R_6_c55, R_6_c56 :  std_logic_vector(2 downto 0);
signal Cin_7_c40, Cin_7_c41 :  std_logic;
signal X_7_c33, X_7_c34, X_7_c35, X_7_c36, X_7_c37, X_7_c38, X_7_c39, X_7_c40, X_7_c41 :  std_logic_vector(3 downto 0);
signal Y_7_c0, Y_7_c1, Y_7_c2, Y_7_c3, Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12, Y_7_c13, Y_7_c14, Y_7_c15, Y_7_c16, Y_7_c17, Y_7_c18, Y_7_c19, Y_7_c20, Y_7_c21, Y_7_c22, Y_7_c23, Y_7_c24, Y_7_c25, Y_7_c26, Y_7_c27, Y_7_c28, Y_7_c29, Y_7_c30, Y_7_c31, Y_7_c32, Y_7_c33, Y_7_c34, Y_7_c35, Y_7_c36, Y_7_c37, Y_7_c38, Y_7_c39, Y_7_c40, Y_7_c41 :  std_logic_vector(3 downto 0);
signal S_7_c41 :  std_logic_vector(3 downto 0);
signal R_7_c41, R_7_c42, R_7_c43, R_7_c44, R_7_c45, R_7_c46, R_7_c47, R_7_c48, R_7_c49, R_7_c50, R_7_c51, R_7_c52, R_7_c53, R_7_c54, R_7_c55, R_7_c56 :  std_logic_vector(2 downto 0);
signal Cin_8_c41, Cin_8_c42 :  std_logic;
signal X_8_c33, X_8_c34, X_8_c35, X_8_c36, X_8_c37, X_8_c38, X_8_c39, X_8_c40, X_8_c41, X_8_c42 :  std_logic_vector(3 downto 0);
signal Y_8_c0, Y_8_c1, Y_8_c2, Y_8_c3, Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13, Y_8_c14, Y_8_c15, Y_8_c16, Y_8_c17, Y_8_c18, Y_8_c19, Y_8_c20, Y_8_c21, Y_8_c22, Y_8_c23, Y_8_c24, Y_8_c25, Y_8_c26, Y_8_c27, Y_8_c28, Y_8_c29, Y_8_c30, Y_8_c31, Y_8_c32, Y_8_c33, Y_8_c34, Y_8_c35, Y_8_c36, Y_8_c37, Y_8_c38, Y_8_c39, Y_8_c40, Y_8_c41, Y_8_c42 :  std_logic_vector(3 downto 0);
signal S_8_c42 :  std_logic_vector(3 downto 0);
signal R_8_c42, R_8_c43, R_8_c44, R_8_c45, R_8_c46, R_8_c47, R_8_c48, R_8_c49, R_8_c50, R_8_c51, R_8_c52, R_8_c53, R_8_c54, R_8_c55, R_8_c56 :  std_logic_vector(2 downto 0);
signal Cin_9_c42, Cin_9_c43 :  std_logic;
signal X_9_c33, X_9_c34, X_9_c35, X_9_c36, X_9_c37, X_9_c38, X_9_c39, X_9_c40, X_9_c41, X_9_c42, X_9_c43 :  std_logic_vector(3 downto 0);
signal Y_9_c0, Y_9_c1, Y_9_c2, Y_9_c3, Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14, Y_9_c15, Y_9_c16, Y_9_c17, Y_9_c18, Y_9_c19, Y_9_c20, Y_9_c21, Y_9_c22, Y_9_c23, Y_9_c24, Y_9_c25, Y_9_c26, Y_9_c27, Y_9_c28, Y_9_c29, Y_9_c30, Y_9_c31, Y_9_c32, Y_9_c33, Y_9_c34, Y_9_c35, Y_9_c36, Y_9_c37, Y_9_c38, Y_9_c39, Y_9_c40, Y_9_c41, Y_9_c42, Y_9_c43 :  std_logic_vector(3 downto 0);
signal S_9_c43 :  std_logic_vector(3 downto 0);
signal R_9_c43, R_9_c44, R_9_c45, R_9_c46, R_9_c47, R_9_c48, R_9_c49, R_9_c50, R_9_c51, R_9_c52, R_9_c53, R_9_c54, R_9_c55, R_9_c56 :  std_logic_vector(2 downto 0);
signal Cin_10_c43, Cin_10_c44 :  std_logic;
signal X_10_c33, X_10_c34, X_10_c35, X_10_c36, X_10_c37, X_10_c38, X_10_c39, X_10_c40, X_10_c41, X_10_c42, X_10_c43, X_10_c44 :  std_logic_vector(3 downto 0);
signal Y_10_c0, Y_10_c1, Y_10_c2, Y_10_c3, Y_10_c4, Y_10_c5, Y_10_c6, Y_10_c7, Y_10_c8, Y_10_c9, Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15, Y_10_c16, Y_10_c17, Y_10_c18, Y_10_c19, Y_10_c20, Y_10_c21, Y_10_c22, Y_10_c23, Y_10_c24, Y_10_c25, Y_10_c26, Y_10_c27, Y_10_c28, Y_10_c29, Y_10_c30, Y_10_c31, Y_10_c32, Y_10_c33, Y_10_c34, Y_10_c35, Y_10_c36, Y_10_c37, Y_10_c38, Y_10_c39, Y_10_c40, Y_10_c41, Y_10_c42, Y_10_c43, Y_10_c44 :  std_logic_vector(3 downto 0);
signal S_10_c44 :  std_logic_vector(3 downto 0);
signal R_10_c44, R_10_c45, R_10_c46, R_10_c47, R_10_c48, R_10_c49, R_10_c50, R_10_c51, R_10_c52, R_10_c53, R_10_c54, R_10_c55, R_10_c56 :  std_logic_vector(2 downto 0);
signal Cin_11_c44, Cin_11_c45 :  std_logic;
signal X_11_c33, X_11_c34, X_11_c35, X_11_c36, X_11_c37, X_11_c38, X_11_c39, X_11_c40, X_11_c41, X_11_c42, X_11_c43, X_11_c44, X_11_c45 :  std_logic_vector(3 downto 0);
signal Y_11_c0, Y_11_c1, Y_11_c2, Y_11_c3, Y_11_c4, Y_11_c5, Y_11_c6, Y_11_c7, Y_11_c8, Y_11_c9, Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16, Y_11_c17, Y_11_c18, Y_11_c19, Y_11_c20, Y_11_c21, Y_11_c22, Y_11_c23, Y_11_c24, Y_11_c25, Y_11_c26, Y_11_c27, Y_11_c28, Y_11_c29, Y_11_c30, Y_11_c31, Y_11_c32, Y_11_c33, Y_11_c34, Y_11_c35, Y_11_c36, Y_11_c37, Y_11_c38, Y_11_c39, Y_11_c40, Y_11_c41, Y_11_c42, Y_11_c43, Y_11_c44, Y_11_c45 :  std_logic_vector(3 downto 0);
signal S_11_c45 :  std_logic_vector(3 downto 0);
signal R_11_c45, R_11_c46, R_11_c47, R_11_c48, R_11_c49, R_11_c50, R_11_c51, R_11_c52, R_11_c53, R_11_c54, R_11_c55, R_11_c56 :  std_logic_vector(2 downto 0);
signal Cin_12_c45, Cin_12_c46 :  std_logic;
signal X_12_c33, X_12_c34, X_12_c35, X_12_c36, X_12_c37, X_12_c38, X_12_c39, X_12_c40, X_12_c41, X_12_c42, X_12_c43, X_12_c44, X_12_c45, X_12_c46 :  std_logic_vector(3 downto 0);
signal Y_12_c0, Y_12_c1, Y_12_c2, Y_12_c3, Y_12_c4, Y_12_c5, Y_12_c6, Y_12_c7, Y_12_c8, Y_12_c9, Y_12_c10, Y_12_c11, Y_12_c12, Y_12_c13, Y_12_c14, Y_12_c15, Y_12_c16, Y_12_c17, Y_12_c18, Y_12_c19, Y_12_c20, Y_12_c21, Y_12_c22, Y_12_c23, Y_12_c24, Y_12_c25, Y_12_c26, Y_12_c27, Y_12_c28, Y_12_c29, Y_12_c30, Y_12_c31, Y_12_c32, Y_12_c33, Y_12_c34, Y_12_c35, Y_12_c36, Y_12_c37, Y_12_c38, Y_12_c39, Y_12_c40, Y_12_c41, Y_12_c42, Y_12_c43, Y_12_c44, Y_12_c45, Y_12_c46 :  std_logic_vector(3 downto 0);
signal S_12_c46 :  std_logic_vector(3 downto 0);
signal R_12_c46, R_12_c47, R_12_c48, R_12_c49, R_12_c50, R_12_c51, R_12_c52, R_12_c53, R_12_c54, R_12_c55, R_12_c56 :  std_logic_vector(2 downto 0);
signal Cin_13_c46, Cin_13_c47 :  std_logic;
signal X_13_c33, X_13_c34, X_13_c35, X_13_c36, X_13_c37, X_13_c38, X_13_c39, X_13_c40, X_13_c41, X_13_c42, X_13_c43, X_13_c44, X_13_c45, X_13_c46, X_13_c47 :  std_logic_vector(3 downto 0);
signal Y_13_c0, Y_13_c1, Y_13_c2, Y_13_c3, Y_13_c4, Y_13_c5, Y_13_c6, Y_13_c7, Y_13_c8, Y_13_c9, Y_13_c10, Y_13_c11, Y_13_c12, Y_13_c13, Y_13_c14, Y_13_c15, Y_13_c16, Y_13_c17, Y_13_c18, Y_13_c19, Y_13_c20, Y_13_c21, Y_13_c22, Y_13_c23, Y_13_c24, Y_13_c25, Y_13_c26, Y_13_c27, Y_13_c28, Y_13_c29, Y_13_c30, Y_13_c31, Y_13_c32, Y_13_c33, Y_13_c34, Y_13_c35, Y_13_c36, Y_13_c37, Y_13_c38, Y_13_c39, Y_13_c40, Y_13_c41, Y_13_c42, Y_13_c43, Y_13_c44, Y_13_c45, Y_13_c46, Y_13_c47 :  std_logic_vector(3 downto 0);
signal S_13_c47 :  std_logic_vector(3 downto 0);
signal R_13_c47, R_13_c48, R_13_c49, R_13_c50, R_13_c51, R_13_c52, R_13_c53, R_13_c54, R_13_c55, R_13_c56 :  std_logic_vector(2 downto 0);
signal Cin_14_c47, Cin_14_c48 :  std_logic;
signal X_14_c33, X_14_c34, X_14_c35, X_14_c36, X_14_c37, X_14_c38, X_14_c39, X_14_c40, X_14_c41, X_14_c42, X_14_c43, X_14_c44, X_14_c45, X_14_c46, X_14_c47, X_14_c48 :  std_logic_vector(3 downto 0);
signal Y_14_c0, Y_14_c1, Y_14_c2, Y_14_c3, Y_14_c4, Y_14_c5, Y_14_c6, Y_14_c7, Y_14_c8, Y_14_c9, Y_14_c10, Y_14_c11, Y_14_c12, Y_14_c13, Y_14_c14, Y_14_c15, Y_14_c16, Y_14_c17, Y_14_c18, Y_14_c19, Y_14_c20, Y_14_c21, Y_14_c22, Y_14_c23, Y_14_c24, Y_14_c25, Y_14_c26, Y_14_c27, Y_14_c28, Y_14_c29, Y_14_c30, Y_14_c31, Y_14_c32, Y_14_c33, Y_14_c34, Y_14_c35, Y_14_c36, Y_14_c37, Y_14_c38, Y_14_c39, Y_14_c40, Y_14_c41, Y_14_c42, Y_14_c43, Y_14_c44, Y_14_c45, Y_14_c46, Y_14_c47, Y_14_c48 :  std_logic_vector(3 downto 0);
signal S_14_c48 :  std_logic_vector(3 downto 0);
signal R_14_c48, R_14_c49, R_14_c50, R_14_c51, R_14_c52, R_14_c53, R_14_c54, R_14_c55, R_14_c56 :  std_logic_vector(2 downto 0);
signal Cin_15_c48, Cin_15_c49 :  std_logic;
signal X_15_c33, X_15_c34, X_15_c35, X_15_c36, X_15_c37, X_15_c38, X_15_c39, X_15_c40, X_15_c41, X_15_c42, X_15_c43, X_15_c44, X_15_c45, X_15_c46, X_15_c47, X_15_c48, X_15_c49 :  std_logic_vector(3 downto 0);
signal Y_15_c0, Y_15_c1, Y_15_c2, Y_15_c3, Y_15_c4, Y_15_c5, Y_15_c6, Y_15_c7, Y_15_c8, Y_15_c9, Y_15_c10, Y_15_c11, Y_15_c12, Y_15_c13, Y_15_c14, Y_15_c15, Y_15_c16, Y_15_c17, Y_15_c18, Y_15_c19, Y_15_c20, Y_15_c21, Y_15_c22, Y_15_c23, Y_15_c24, Y_15_c25, Y_15_c26, Y_15_c27, Y_15_c28, Y_15_c29, Y_15_c30, Y_15_c31, Y_15_c32, Y_15_c33, Y_15_c34, Y_15_c35, Y_15_c36, Y_15_c37, Y_15_c38, Y_15_c39, Y_15_c40, Y_15_c41, Y_15_c42, Y_15_c43, Y_15_c44, Y_15_c45, Y_15_c46, Y_15_c47, Y_15_c48, Y_15_c49 :  std_logic_vector(3 downto 0);
signal S_15_c49 :  std_logic_vector(3 downto 0);
signal R_15_c49, R_15_c50, R_15_c51, R_15_c52, R_15_c53, R_15_c54, R_15_c55, R_15_c56 :  std_logic_vector(2 downto 0);
signal Cin_16_c49, Cin_16_c50 :  std_logic;
signal X_16_c33, X_16_c34, X_16_c35, X_16_c36, X_16_c37, X_16_c38, X_16_c39, X_16_c40, X_16_c41, X_16_c42, X_16_c43, X_16_c44, X_16_c45, X_16_c46, X_16_c47, X_16_c48, X_16_c49, X_16_c50 :  std_logic_vector(3 downto 0);
signal Y_16_c0, Y_16_c1, Y_16_c2, Y_16_c3, Y_16_c4, Y_16_c5, Y_16_c6, Y_16_c7, Y_16_c8, Y_16_c9, Y_16_c10, Y_16_c11, Y_16_c12, Y_16_c13, Y_16_c14, Y_16_c15, Y_16_c16, Y_16_c17, Y_16_c18, Y_16_c19, Y_16_c20, Y_16_c21, Y_16_c22, Y_16_c23, Y_16_c24, Y_16_c25, Y_16_c26, Y_16_c27, Y_16_c28, Y_16_c29, Y_16_c30, Y_16_c31, Y_16_c32, Y_16_c33, Y_16_c34, Y_16_c35, Y_16_c36, Y_16_c37, Y_16_c38, Y_16_c39, Y_16_c40, Y_16_c41, Y_16_c42, Y_16_c43, Y_16_c44, Y_16_c45, Y_16_c46, Y_16_c47, Y_16_c48, Y_16_c49, Y_16_c50 :  std_logic_vector(3 downto 0);
signal S_16_c50 :  std_logic_vector(3 downto 0);
signal R_16_c50, R_16_c51, R_16_c52, R_16_c53, R_16_c54, R_16_c55, R_16_c56 :  std_logic_vector(2 downto 0);
signal Cin_17_c50, Cin_17_c51 :  std_logic;
signal X_17_c33, X_17_c34, X_17_c35, X_17_c36, X_17_c37, X_17_c38, X_17_c39, X_17_c40, X_17_c41, X_17_c42, X_17_c43, X_17_c44, X_17_c45, X_17_c46, X_17_c47, X_17_c48, X_17_c49, X_17_c50, X_17_c51 :  std_logic_vector(3 downto 0);
signal Y_17_c0, Y_17_c1, Y_17_c2, Y_17_c3, Y_17_c4, Y_17_c5, Y_17_c6, Y_17_c7, Y_17_c8, Y_17_c9, Y_17_c10, Y_17_c11, Y_17_c12, Y_17_c13, Y_17_c14, Y_17_c15, Y_17_c16, Y_17_c17, Y_17_c18, Y_17_c19, Y_17_c20, Y_17_c21, Y_17_c22, Y_17_c23, Y_17_c24, Y_17_c25, Y_17_c26, Y_17_c27, Y_17_c28, Y_17_c29, Y_17_c30, Y_17_c31, Y_17_c32, Y_17_c33, Y_17_c34, Y_17_c35, Y_17_c36, Y_17_c37, Y_17_c38, Y_17_c39, Y_17_c40, Y_17_c41, Y_17_c42, Y_17_c43, Y_17_c44, Y_17_c45, Y_17_c46, Y_17_c47, Y_17_c48, Y_17_c49, Y_17_c50, Y_17_c51 :  std_logic_vector(3 downto 0);
signal S_17_c51 :  std_logic_vector(3 downto 0);
signal R_17_c51, R_17_c52, R_17_c53, R_17_c54, R_17_c55, R_17_c56 :  std_logic_vector(2 downto 0);
signal Cin_18_c51, Cin_18_c52 :  std_logic;
signal X_18_c33, X_18_c34, X_18_c35, X_18_c36, X_18_c37, X_18_c38, X_18_c39, X_18_c40, X_18_c41, X_18_c42, X_18_c43, X_18_c44, X_18_c45, X_18_c46, X_18_c47, X_18_c48, X_18_c49, X_18_c50, X_18_c51, X_18_c52 :  std_logic_vector(3 downto 0);
signal Y_18_c0, Y_18_c1, Y_18_c2, Y_18_c3, Y_18_c4, Y_18_c5, Y_18_c6, Y_18_c7, Y_18_c8, Y_18_c9, Y_18_c10, Y_18_c11, Y_18_c12, Y_18_c13, Y_18_c14, Y_18_c15, Y_18_c16, Y_18_c17, Y_18_c18, Y_18_c19, Y_18_c20, Y_18_c21, Y_18_c22, Y_18_c23, Y_18_c24, Y_18_c25, Y_18_c26, Y_18_c27, Y_18_c28, Y_18_c29, Y_18_c30, Y_18_c31, Y_18_c32, Y_18_c33, Y_18_c34, Y_18_c35, Y_18_c36, Y_18_c37, Y_18_c38, Y_18_c39, Y_18_c40, Y_18_c41, Y_18_c42, Y_18_c43, Y_18_c44, Y_18_c45, Y_18_c46, Y_18_c47, Y_18_c48, Y_18_c49, Y_18_c50, Y_18_c51, Y_18_c52 :  std_logic_vector(3 downto 0);
signal S_18_c52 :  std_logic_vector(3 downto 0);
signal R_18_c52, R_18_c53, R_18_c54, R_18_c55, R_18_c56 :  std_logic_vector(2 downto 0);
signal Cin_19_c52, Cin_19_c53 :  std_logic;
signal X_19_c33, X_19_c34, X_19_c35, X_19_c36, X_19_c37, X_19_c38, X_19_c39, X_19_c40, X_19_c41, X_19_c42, X_19_c43, X_19_c44, X_19_c45, X_19_c46, X_19_c47, X_19_c48, X_19_c49, X_19_c50, X_19_c51, X_19_c52, X_19_c53 :  std_logic_vector(3 downto 0);
signal Y_19_c0, Y_19_c1, Y_19_c2, Y_19_c3, Y_19_c4, Y_19_c5, Y_19_c6, Y_19_c7, Y_19_c8, Y_19_c9, Y_19_c10, Y_19_c11, Y_19_c12, Y_19_c13, Y_19_c14, Y_19_c15, Y_19_c16, Y_19_c17, Y_19_c18, Y_19_c19, Y_19_c20, Y_19_c21, Y_19_c22, Y_19_c23, Y_19_c24, Y_19_c25, Y_19_c26, Y_19_c27, Y_19_c28, Y_19_c29, Y_19_c30, Y_19_c31, Y_19_c32, Y_19_c33, Y_19_c34, Y_19_c35, Y_19_c36, Y_19_c37, Y_19_c38, Y_19_c39, Y_19_c40, Y_19_c41, Y_19_c42, Y_19_c43, Y_19_c44, Y_19_c45, Y_19_c46, Y_19_c47, Y_19_c48, Y_19_c49, Y_19_c50, Y_19_c51, Y_19_c52, Y_19_c53 :  std_logic_vector(3 downto 0);
signal S_19_c53 :  std_logic_vector(3 downto 0);
signal R_19_c53, R_19_c54, R_19_c55, R_19_c56 :  std_logic_vector(2 downto 0);
signal Cin_20_c53, Cin_20_c54 :  std_logic;
signal X_20_c33, X_20_c34, X_20_c35, X_20_c36, X_20_c37, X_20_c38, X_20_c39, X_20_c40, X_20_c41, X_20_c42, X_20_c43, X_20_c44, X_20_c45, X_20_c46, X_20_c47, X_20_c48, X_20_c49, X_20_c50, X_20_c51, X_20_c52, X_20_c53, X_20_c54 :  std_logic_vector(3 downto 0);
signal Y_20_c0, Y_20_c1, Y_20_c2, Y_20_c3, Y_20_c4, Y_20_c5, Y_20_c6, Y_20_c7, Y_20_c8, Y_20_c9, Y_20_c10, Y_20_c11, Y_20_c12, Y_20_c13, Y_20_c14, Y_20_c15, Y_20_c16, Y_20_c17, Y_20_c18, Y_20_c19, Y_20_c20, Y_20_c21, Y_20_c22, Y_20_c23, Y_20_c24, Y_20_c25, Y_20_c26, Y_20_c27, Y_20_c28, Y_20_c29, Y_20_c30, Y_20_c31, Y_20_c32, Y_20_c33, Y_20_c34, Y_20_c35, Y_20_c36, Y_20_c37, Y_20_c38, Y_20_c39, Y_20_c40, Y_20_c41, Y_20_c42, Y_20_c43, Y_20_c44, Y_20_c45, Y_20_c46, Y_20_c47, Y_20_c48, Y_20_c49, Y_20_c50, Y_20_c51, Y_20_c52, Y_20_c53, Y_20_c54 :  std_logic_vector(3 downto 0);
signal S_20_c54 :  std_logic_vector(3 downto 0);
signal R_20_c54, R_20_c55, R_20_c56 :  std_logic_vector(2 downto 0);
signal Cin_21_c54, Cin_21_c55, Cin_21_c56 :  std_logic;
signal X_21_c33, X_21_c34, X_21_c35, X_21_c36, X_21_c37, X_21_c38, X_21_c39, X_21_c40, X_21_c41, X_21_c42, X_21_c43, X_21_c44, X_21_c45, X_21_c46, X_21_c47, X_21_c48, X_21_c49, X_21_c50, X_21_c51, X_21_c52, X_21_c53, X_21_c54, X_21_c55, X_21_c56 :  std_logic_vector(3 downto 0);
signal Y_21_c0, Y_21_c1, Y_21_c2, Y_21_c3, Y_21_c4, Y_21_c5, Y_21_c6, Y_21_c7, Y_21_c8, Y_21_c9, Y_21_c10, Y_21_c11, Y_21_c12, Y_21_c13, Y_21_c14, Y_21_c15, Y_21_c16, Y_21_c17, Y_21_c18, Y_21_c19, Y_21_c20, Y_21_c21, Y_21_c22, Y_21_c23, Y_21_c24, Y_21_c25, Y_21_c26, Y_21_c27, Y_21_c28, Y_21_c29, Y_21_c30, Y_21_c31, Y_21_c32, Y_21_c33, Y_21_c34, Y_21_c35, Y_21_c36, Y_21_c37, Y_21_c38, Y_21_c39, Y_21_c40, Y_21_c41, Y_21_c42, Y_21_c43, Y_21_c44, Y_21_c45, Y_21_c46, Y_21_c47, Y_21_c48, Y_21_c49, Y_21_c50, Y_21_c51, Y_21_c52, Y_21_c53, Y_21_c54, Y_21_c55, Y_21_c56 :  std_logic_vector(3 downto 0);
signal S_21_c56 :  std_logic_vector(3 downto 0);
signal R_21_c56 :  std_logic_vector(2 downto 0);
signal Cin_22_c56 :  std_logic;
signal X_22_c33, X_22_c34, X_22_c35, X_22_c36, X_22_c37, X_22_c38, X_22_c39, X_22_c40, X_22_c41, X_22_c42, X_22_c43, X_22_c44, X_22_c45, X_22_c46, X_22_c47, X_22_c48, X_22_c49, X_22_c50, X_22_c51, X_22_c52, X_22_c53, X_22_c54, X_22_c55, X_22_c56 :  std_logic_vector(2 downto 0);
signal Y_22_c0, Y_22_c1, Y_22_c2, Y_22_c3, Y_22_c4, Y_22_c5, Y_22_c6, Y_22_c7, Y_22_c8, Y_22_c9, Y_22_c10, Y_22_c11, Y_22_c12, Y_22_c13, Y_22_c14, Y_22_c15, Y_22_c16, Y_22_c17, Y_22_c18, Y_22_c19, Y_22_c20, Y_22_c21, Y_22_c22, Y_22_c23, Y_22_c24, Y_22_c25, Y_22_c26, Y_22_c27, Y_22_c28, Y_22_c29, Y_22_c30, Y_22_c31, Y_22_c32, Y_22_c33, Y_22_c34, Y_22_c35, Y_22_c36, Y_22_c37, Y_22_c38, Y_22_c39, Y_22_c40, Y_22_c41, Y_22_c42, Y_22_c43, Y_22_c44, Y_22_c45, Y_22_c46, Y_22_c47, Y_22_c48, Y_22_c49, Y_22_c50, Y_22_c51, Y_22_c52, Y_22_c53, Y_22_c54, Y_22_c55, Y_22_c56 :  std_logic_vector(2 downto 0);
signal S_22_c56 :  std_logic_vector(2 downto 0);
signal R_22_c56 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
               Y_2_c1 <= Y_2_c0;
               Y_3_c1 <= Y_3_c0;
               Y_4_c1 <= Y_4_c0;
               Y_5_c1 <= Y_5_c0;
               Y_6_c1 <= Y_6_c0;
               Y_7_c1 <= Y_7_c0;
               Y_8_c1 <= Y_8_c0;
               Y_9_c1 <= Y_9_c0;
               Y_10_c1 <= Y_10_c0;
               Y_11_c1 <= Y_11_c0;
               Y_12_c1 <= Y_12_c0;
               Y_13_c1 <= Y_13_c0;
               Y_14_c1 <= Y_14_c0;
               Y_15_c1 <= Y_15_c0;
               Y_16_c1 <= Y_16_c0;
               Y_17_c1 <= Y_17_c0;
               Y_18_c1 <= Y_18_c0;
               Y_19_c1 <= Y_19_c0;
               Y_20_c1 <= Y_20_c0;
               Y_21_c1 <= Y_21_c0;
               Y_22_c1 <= Y_22_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
               Y_2_c2 <= Y_2_c1;
               Y_3_c2 <= Y_3_c1;
               Y_4_c2 <= Y_4_c1;
               Y_5_c2 <= Y_5_c1;
               Y_6_c2 <= Y_6_c1;
               Y_7_c2 <= Y_7_c1;
               Y_8_c2 <= Y_8_c1;
               Y_9_c2 <= Y_9_c1;
               Y_10_c2 <= Y_10_c1;
               Y_11_c2 <= Y_11_c1;
               Y_12_c2 <= Y_12_c1;
               Y_13_c2 <= Y_13_c1;
               Y_14_c2 <= Y_14_c1;
               Y_15_c2 <= Y_15_c1;
               Y_16_c2 <= Y_16_c1;
               Y_17_c2 <= Y_17_c1;
               Y_18_c2 <= Y_18_c1;
               Y_19_c2 <= Y_19_c1;
               Y_20_c2 <= Y_20_c1;
               Y_21_c2 <= Y_21_c1;
               Y_22_c2 <= Y_22_c1;
            end if;
            if ce_3 = '1' then
               Y_1_c3 <= Y_1_c2;
               Y_2_c3 <= Y_2_c2;
               Y_3_c3 <= Y_3_c2;
               Y_4_c3 <= Y_4_c2;
               Y_5_c3 <= Y_5_c2;
               Y_6_c3 <= Y_6_c2;
               Y_7_c3 <= Y_7_c2;
               Y_8_c3 <= Y_8_c2;
               Y_9_c3 <= Y_9_c2;
               Y_10_c3 <= Y_10_c2;
               Y_11_c3 <= Y_11_c2;
               Y_12_c3 <= Y_12_c2;
               Y_13_c3 <= Y_13_c2;
               Y_14_c3 <= Y_14_c2;
               Y_15_c3 <= Y_15_c2;
               Y_16_c3 <= Y_16_c2;
               Y_17_c3 <= Y_17_c2;
               Y_18_c3 <= Y_18_c2;
               Y_19_c3 <= Y_19_c2;
               Y_20_c3 <= Y_20_c2;
               Y_21_c3 <= Y_21_c2;
               Y_22_c3 <= Y_22_c2;
            end if;
            if ce_4 = '1' then
               Y_1_c4 <= Y_1_c3;
               Y_2_c4 <= Y_2_c3;
               Y_3_c4 <= Y_3_c3;
               Y_4_c4 <= Y_4_c3;
               Y_5_c4 <= Y_5_c3;
               Y_6_c4 <= Y_6_c3;
               Y_7_c4 <= Y_7_c3;
               Y_8_c4 <= Y_8_c3;
               Y_9_c4 <= Y_9_c3;
               Y_10_c4 <= Y_10_c3;
               Y_11_c4 <= Y_11_c3;
               Y_12_c4 <= Y_12_c3;
               Y_13_c4 <= Y_13_c3;
               Y_14_c4 <= Y_14_c3;
               Y_15_c4 <= Y_15_c3;
               Y_16_c4 <= Y_16_c3;
               Y_17_c4 <= Y_17_c3;
               Y_18_c4 <= Y_18_c3;
               Y_19_c4 <= Y_19_c3;
               Y_20_c4 <= Y_20_c3;
               Y_21_c4 <= Y_21_c3;
               Y_22_c4 <= Y_22_c3;
            end if;
            if ce_5 = '1' then
               Y_1_c5 <= Y_1_c4;
               Y_2_c5 <= Y_2_c4;
               Y_3_c5 <= Y_3_c4;
               Y_4_c5 <= Y_4_c4;
               Y_5_c5 <= Y_5_c4;
               Y_6_c5 <= Y_6_c4;
               Y_7_c5 <= Y_7_c4;
               Y_8_c5 <= Y_8_c4;
               Y_9_c5 <= Y_9_c4;
               Y_10_c5 <= Y_10_c4;
               Y_11_c5 <= Y_11_c4;
               Y_12_c5 <= Y_12_c4;
               Y_13_c5 <= Y_13_c4;
               Y_14_c5 <= Y_14_c4;
               Y_15_c5 <= Y_15_c4;
               Y_16_c5 <= Y_16_c4;
               Y_17_c5 <= Y_17_c4;
               Y_18_c5 <= Y_18_c4;
               Y_19_c5 <= Y_19_c4;
               Y_20_c5 <= Y_20_c4;
               Y_21_c5 <= Y_21_c4;
               Y_22_c5 <= Y_22_c4;
            end if;
            if ce_6 = '1' then
               Y_1_c6 <= Y_1_c5;
               Y_2_c6 <= Y_2_c5;
               Y_3_c6 <= Y_3_c5;
               Y_4_c6 <= Y_4_c5;
               Y_5_c6 <= Y_5_c5;
               Y_6_c6 <= Y_6_c5;
               Y_7_c6 <= Y_7_c5;
               Y_8_c6 <= Y_8_c5;
               Y_9_c6 <= Y_9_c5;
               Y_10_c6 <= Y_10_c5;
               Y_11_c6 <= Y_11_c5;
               Y_12_c6 <= Y_12_c5;
               Y_13_c6 <= Y_13_c5;
               Y_14_c6 <= Y_14_c5;
               Y_15_c6 <= Y_15_c5;
               Y_16_c6 <= Y_16_c5;
               Y_17_c6 <= Y_17_c5;
               Y_18_c6 <= Y_18_c5;
               Y_19_c6 <= Y_19_c5;
               Y_20_c6 <= Y_20_c5;
               Y_21_c6 <= Y_21_c5;
               Y_22_c6 <= Y_22_c5;
            end if;
            if ce_7 = '1' then
               Y_1_c7 <= Y_1_c6;
               Y_2_c7 <= Y_2_c6;
               Y_3_c7 <= Y_3_c6;
               Y_4_c7 <= Y_4_c6;
               Y_5_c7 <= Y_5_c6;
               Y_6_c7 <= Y_6_c6;
               Y_7_c7 <= Y_7_c6;
               Y_8_c7 <= Y_8_c6;
               Y_9_c7 <= Y_9_c6;
               Y_10_c7 <= Y_10_c6;
               Y_11_c7 <= Y_11_c6;
               Y_12_c7 <= Y_12_c6;
               Y_13_c7 <= Y_13_c6;
               Y_14_c7 <= Y_14_c6;
               Y_15_c7 <= Y_15_c6;
               Y_16_c7 <= Y_16_c6;
               Y_17_c7 <= Y_17_c6;
               Y_18_c7 <= Y_18_c6;
               Y_19_c7 <= Y_19_c6;
               Y_20_c7 <= Y_20_c6;
               Y_21_c7 <= Y_21_c6;
               Y_22_c7 <= Y_22_c6;
            end if;
            if ce_8 = '1' then
               Y_1_c8 <= Y_1_c7;
               Y_2_c8 <= Y_2_c7;
               Y_3_c8 <= Y_3_c7;
               Y_4_c8 <= Y_4_c7;
               Y_5_c8 <= Y_5_c7;
               Y_6_c8 <= Y_6_c7;
               Y_7_c8 <= Y_7_c7;
               Y_8_c8 <= Y_8_c7;
               Y_9_c8 <= Y_9_c7;
               Y_10_c8 <= Y_10_c7;
               Y_11_c8 <= Y_11_c7;
               Y_12_c8 <= Y_12_c7;
               Y_13_c8 <= Y_13_c7;
               Y_14_c8 <= Y_14_c7;
               Y_15_c8 <= Y_15_c7;
               Y_16_c8 <= Y_16_c7;
               Y_17_c8 <= Y_17_c7;
               Y_18_c8 <= Y_18_c7;
               Y_19_c8 <= Y_19_c7;
               Y_20_c8 <= Y_20_c7;
               Y_21_c8 <= Y_21_c7;
               Y_22_c8 <= Y_22_c7;
            end if;
            if ce_9 = '1' then
               Y_1_c9 <= Y_1_c8;
               Y_2_c9 <= Y_2_c8;
               Y_3_c9 <= Y_3_c8;
               Y_4_c9 <= Y_4_c8;
               Y_5_c9 <= Y_5_c8;
               Y_6_c9 <= Y_6_c8;
               Y_7_c9 <= Y_7_c8;
               Y_8_c9 <= Y_8_c8;
               Y_9_c9 <= Y_9_c8;
               Y_10_c9 <= Y_10_c8;
               Y_11_c9 <= Y_11_c8;
               Y_12_c9 <= Y_12_c8;
               Y_13_c9 <= Y_13_c8;
               Y_14_c9 <= Y_14_c8;
               Y_15_c9 <= Y_15_c8;
               Y_16_c9 <= Y_16_c8;
               Y_17_c9 <= Y_17_c8;
               Y_18_c9 <= Y_18_c8;
               Y_19_c9 <= Y_19_c8;
               Y_20_c9 <= Y_20_c8;
               Y_21_c9 <= Y_21_c8;
               Y_22_c9 <= Y_22_c8;
            end if;
            if ce_10 = '1' then
               Y_1_c10 <= Y_1_c9;
               Y_2_c10 <= Y_2_c9;
               Y_3_c10 <= Y_3_c9;
               Y_4_c10 <= Y_4_c9;
               Y_5_c10 <= Y_5_c9;
               Y_6_c10 <= Y_6_c9;
               Y_7_c10 <= Y_7_c9;
               Y_8_c10 <= Y_8_c9;
               Y_9_c10 <= Y_9_c9;
               Y_10_c10 <= Y_10_c9;
               Y_11_c10 <= Y_11_c9;
               Y_12_c10 <= Y_12_c9;
               Y_13_c10 <= Y_13_c9;
               Y_14_c10 <= Y_14_c9;
               Y_15_c10 <= Y_15_c9;
               Y_16_c10 <= Y_16_c9;
               Y_17_c10 <= Y_17_c9;
               Y_18_c10 <= Y_18_c9;
               Y_19_c10 <= Y_19_c9;
               Y_20_c10 <= Y_20_c9;
               Y_21_c10 <= Y_21_c9;
               Y_22_c10 <= Y_22_c9;
            end if;
            if ce_11 = '1' then
               Y_1_c11 <= Y_1_c10;
               Y_2_c11 <= Y_2_c10;
               Y_3_c11 <= Y_3_c10;
               Y_4_c11 <= Y_4_c10;
               Y_5_c11 <= Y_5_c10;
               Y_6_c11 <= Y_6_c10;
               Y_7_c11 <= Y_7_c10;
               Y_8_c11 <= Y_8_c10;
               Y_9_c11 <= Y_9_c10;
               Y_10_c11 <= Y_10_c10;
               Y_11_c11 <= Y_11_c10;
               Y_12_c11 <= Y_12_c10;
               Y_13_c11 <= Y_13_c10;
               Y_14_c11 <= Y_14_c10;
               Y_15_c11 <= Y_15_c10;
               Y_16_c11 <= Y_16_c10;
               Y_17_c11 <= Y_17_c10;
               Y_18_c11 <= Y_18_c10;
               Y_19_c11 <= Y_19_c10;
               Y_20_c11 <= Y_20_c10;
               Y_21_c11 <= Y_21_c10;
               Y_22_c11 <= Y_22_c10;
            end if;
            if ce_12 = '1' then
               Y_1_c12 <= Y_1_c11;
               Y_2_c12 <= Y_2_c11;
               Y_3_c12 <= Y_3_c11;
               Y_4_c12 <= Y_4_c11;
               Y_5_c12 <= Y_5_c11;
               Y_6_c12 <= Y_6_c11;
               Y_7_c12 <= Y_7_c11;
               Y_8_c12 <= Y_8_c11;
               Y_9_c12 <= Y_9_c11;
               Y_10_c12 <= Y_10_c11;
               Y_11_c12 <= Y_11_c11;
               Y_12_c12 <= Y_12_c11;
               Y_13_c12 <= Y_13_c11;
               Y_14_c12 <= Y_14_c11;
               Y_15_c12 <= Y_15_c11;
               Y_16_c12 <= Y_16_c11;
               Y_17_c12 <= Y_17_c11;
               Y_18_c12 <= Y_18_c11;
               Y_19_c12 <= Y_19_c11;
               Y_20_c12 <= Y_20_c11;
               Y_21_c12 <= Y_21_c11;
               Y_22_c12 <= Y_22_c11;
            end if;
            if ce_13 = '1' then
               Y_1_c13 <= Y_1_c12;
               Y_2_c13 <= Y_2_c12;
               Y_3_c13 <= Y_3_c12;
               Y_4_c13 <= Y_4_c12;
               Y_5_c13 <= Y_5_c12;
               Y_6_c13 <= Y_6_c12;
               Y_7_c13 <= Y_7_c12;
               Y_8_c13 <= Y_8_c12;
               Y_9_c13 <= Y_9_c12;
               Y_10_c13 <= Y_10_c12;
               Y_11_c13 <= Y_11_c12;
               Y_12_c13 <= Y_12_c12;
               Y_13_c13 <= Y_13_c12;
               Y_14_c13 <= Y_14_c12;
               Y_15_c13 <= Y_15_c12;
               Y_16_c13 <= Y_16_c12;
               Y_17_c13 <= Y_17_c12;
               Y_18_c13 <= Y_18_c12;
               Y_19_c13 <= Y_19_c12;
               Y_20_c13 <= Y_20_c12;
               Y_21_c13 <= Y_21_c12;
               Y_22_c13 <= Y_22_c12;
            end if;
            if ce_14 = '1' then
               Y_1_c14 <= Y_1_c13;
               Y_2_c14 <= Y_2_c13;
               Y_3_c14 <= Y_3_c13;
               Y_4_c14 <= Y_4_c13;
               Y_5_c14 <= Y_5_c13;
               Y_6_c14 <= Y_6_c13;
               Y_7_c14 <= Y_7_c13;
               Y_8_c14 <= Y_8_c13;
               Y_9_c14 <= Y_9_c13;
               Y_10_c14 <= Y_10_c13;
               Y_11_c14 <= Y_11_c13;
               Y_12_c14 <= Y_12_c13;
               Y_13_c14 <= Y_13_c13;
               Y_14_c14 <= Y_14_c13;
               Y_15_c14 <= Y_15_c13;
               Y_16_c14 <= Y_16_c13;
               Y_17_c14 <= Y_17_c13;
               Y_18_c14 <= Y_18_c13;
               Y_19_c14 <= Y_19_c13;
               Y_20_c14 <= Y_20_c13;
               Y_21_c14 <= Y_21_c13;
               Y_22_c14 <= Y_22_c13;
            end if;
            if ce_15 = '1' then
               Y_1_c15 <= Y_1_c14;
               Y_2_c15 <= Y_2_c14;
               Y_3_c15 <= Y_3_c14;
               Y_4_c15 <= Y_4_c14;
               Y_5_c15 <= Y_5_c14;
               Y_6_c15 <= Y_6_c14;
               Y_7_c15 <= Y_7_c14;
               Y_8_c15 <= Y_8_c14;
               Y_9_c15 <= Y_9_c14;
               Y_10_c15 <= Y_10_c14;
               Y_11_c15 <= Y_11_c14;
               Y_12_c15 <= Y_12_c14;
               Y_13_c15 <= Y_13_c14;
               Y_14_c15 <= Y_14_c14;
               Y_15_c15 <= Y_15_c14;
               Y_16_c15 <= Y_16_c14;
               Y_17_c15 <= Y_17_c14;
               Y_18_c15 <= Y_18_c14;
               Y_19_c15 <= Y_19_c14;
               Y_20_c15 <= Y_20_c14;
               Y_21_c15 <= Y_21_c14;
               Y_22_c15 <= Y_22_c14;
            end if;
            if ce_16 = '1' then
               Y_1_c16 <= Y_1_c15;
               Y_2_c16 <= Y_2_c15;
               Y_3_c16 <= Y_3_c15;
               Y_4_c16 <= Y_4_c15;
               Y_5_c16 <= Y_5_c15;
               Y_6_c16 <= Y_6_c15;
               Y_7_c16 <= Y_7_c15;
               Y_8_c16 <= Y_8_c15;
               Y_9_c16 <= Y_9_c15;
               Y_10_c16 <= Y_10_c15;
               Y_11_c16 <= Y_11_c15;
               Y_12_c16 <= Y_12_c15;
               Y_13_c16 <= Y_13_c15;
               Y_14_c16 <= Y_14_c15;
               Y_15_c16 <= Y_15_c15;
               Y_16_c16 <= Y_16_c15;
               Y_17_c16 <= Y_17_c15;
               Y_18_c16 <= Y_18_c15;
               Y_19_c16 <= Y_19_c15;
               Y_20_c16 <= Y_20_c15;
               Y_21_c16 <= Y_21_c15;
               Y_22_c16 <= Y_22_c15;
            end if;
            if ce_17 = '1' then
               Y_1_c17 <= Y_1_c16;
               Y_2_c17 <= Y_2_c16;
               Y_3_c17 <= Y_3_c16;
               Y_4_c17 <= Y_4_c16;
               Y_5_c17 <= Y_5_c16;
               Y_6_c17 <= Y_6_c16;
               Y_7_c17 <= Y_7_c16;
               Y_8_c17 <= Y_8_c16;
               Y_9_c17 <= Y_9_c16;
               Y_10_c17 <= Y_10_c16;
               Y_11_c17 <= Y_11_c16;
               Y_12_c17 <= Y_12_c16;
               Y_13_c17 <= Y_13_c16;
               Y_14_c17 <= Y_14_c16;
               Y_15_c17 <= Y_15_c16;
               Y_16_c17 <= Y_16_c16;
               Y_17_c17 <= Y_17_c16;
               Y_18_c17 <= Y_18_c16;
               Y_19_c17 <= Y_19_c16;
               Y_20_c17 <= Y_20_c16;
               Y_21_c17 <= Y_21_c16;
               Y_22_c17 <= Y_22_c16;
            end if;
            if ce_18 = '1' then
               Y_1_c18 <= Y_1_c17;
               Y_2_c18 <= Y_2_c17;
               Y_3_c18 <= Y_3_c17;
               Y_4_c18 <= Y_4_c17;
               Y_5_c18 <= Y_5_c17;
               Y_6_c18 <= Y_6_c17;
               Y_7_c18 <= Y_7_c17;
               Y_8_c18 <= Y_8_c17;
               Y_9_c18 <= Y_9_c17;
               Y_10_c18 <= Y_10_c17;
               Y_11_c18 <= Y_11_c17;
               Y_12_c18 <= Y_12_c17;
               Y_13_c18 <= Y_13_c17;
               Y_14_c18 <= Y_14_c17;
               Y_15_c18 <= Y_15_c17;
               Y_16_c18 <= Y_16_c17;
               Y_17_c18 <= Y_17_c17;
               Y_18_c18 <= Y_18_c17;
               Y_19_c18 <= Y_19_c17;
               Y_20_c18 <= Y_20_c17;
               Y_21_c18 <= Y_21_c17;
               Y_22_c18 <= Y_22_c17;
            end if;
            if ce_19 = '1' then
               Y_1_c19 <= Y_1_c18;
               Y_2_c19 <= Y_2_c18;
               Y_3_c19 <= Y_3_c18;
               Y_4_c19 <= Y_4_c18;
               Y_5_c19 <= Y_5_c18;
               Y_6_c19 <= Y_6_c18;
               Y_7_c19 <= Y_7_c18;
               Y_8_c19 <= Y_8_c18;
               Y_9_c19 <= Y_9_c18;
               Y_10_c19 <= Y_10_c18;
               Y_11_c19 <= Y_11_c18;
               Y_12_c19 <= Y_12_c18;
               Y_13_c19 <= Y_13_c18;
               Y_14_c19 <= Y_14_c18;
               Y_15_c19 <= Y_15_c18;
               Y_16_c19 <= Y_16_c18;
               Y_17_c19 <= Y_17_c18;
               Y_18_c19 <= Y_18_c18;
               Y_19_c19 <= Y_19_c18;
               Y_20_c19 <= Y_20_c18;
               Y_21_c19 <= Y_21_c18;
               Y_22_c19 <= Y_22_c18;
            end if;
            if ce_20 = '1' then
               Y_1_c20 <= Y_1_c19;
               Y_2_c20 <= Y_2_c19;
               Y_3_c20 <= Y_3_c19;
               Y_4_c20 <= Y_4_c19;
               Y_5_c20 <= Y_5_c19;
               Y_6_c20 <= Y_6_c19;
               Y_7_c20 <= Y_7_c19;
               Y_8_c20 <= Y_8_c19;
               Y_9_c20 <= Y_9_c19;
               Y_10_c20 <= Y_10_c19;
               Y_11_c20 <= Y_11_c19;
               Y_12_c20 <= Y_12_c19;
               Y_13_c20 <= Y_13_c19;
               Y_14_c20 <= Y_14_c19;
               Y_15_c20 <= Y_15_c19;
               Y_16_c20 <= Y_16_c19;
               Y_17_c20 <= Y_17_c19;
               Y_18_c20 <= Y_18_c19;
               Y_19_c20 <= Y_19_c19;
               Y_20_c20 <= Y_20_c19;
               Y_21_c20 <= Y_21_c19;
               Y_22_c20 <= Y_22_c19;
            end if;
            if ce_21 = '1' then
               Y_1_c21 <= Y_1_c20;
               Y_2_c21 <= Y_2_c20;
               Y_3_c21 <= Y_3_c20;
               Y_4_c21 <= Y_4_c20;
               Y_5_c21 <= Y_5_c20;
               Y_6_c21 <= Y_6_c20;
               Y_7_c21 <= Y_7_c20;
               Y_8_c21 <= Y_8_c20;
               Y_9_c21 <= Y_9_c20;
               Y_10_c21 <= Y_10_c20;
               Y_11_c21 <= Y_11_c20;
               Y_12_c21 <= Y_12_c20;
               Y_13_c21 <= Y_13_c20;
               Y_14_c21 <= Y_14_c20;
               Y_15_c21 <= Y_15_c20;
               Y_16_c21 <= Y_16_c20;
               Y_17_c21 <= Y_17_c20;
               Y_18_c21 <= Y_18_c20;
               Y_19_c21 <= Y_19_c20;
               Y_20_c21 <= Y_20_c20;
               Y_21_c21 <= Y_21_c20;
               Y_22_c21 <= Y_22_c20;
            end if;
            if ce_22 = '1' then
               Y_1_c22 <= Y_1_c21;
               Y_2_c22 <= Y_2_c21;
               Y_3_c22 <= Y_3_c21;
               Y_4_c22 <= Y_4_c21;
               Y_5_c22 <= Y_5_c21;
               Y_6_c22 <= Y_6_c21;
               Y_7_c22 <= Y_7_c21;
               Y_8_c22 <= Y_8_c21;
               Y_9_c22 <= Y_9_c21;
               Y_10_c22 <= Y_10_c21;
               Y_11_c22 <= Y_11_c21;
               Y_12_c22 <= Y_12_c21;
               Y_13_c22 <= Y_13_c21;
               Y_14_c22 <= Y_14_c21;
               Y_15_c22 <= Y_15_c21;
               Y_16_c22 <= Y_16_c21;
               Y_17_c22 <= Y_17_c21;
               Y_18_c22 <= Y_18_c21;
               Y_19_c22 <= Y_19_c21;
               Y_20_c22 <= Y_20_c21;
               Y_21_c22 <= Y_21_c21;
               Y_22_c22 <= Y_22_c21;
            end if;
            if ce_23 = '1' then
               Y_1_c23 <= Y_1_c22;
               Y_2_c23 <= Y_2_c22;
               Y_3_c23 <= Y_3_c22;
               Y_4_c23 <= Y_4_c22;
               Y_5_c23 <= Y_5_c22;
               Y_6_c23 <= Y_6_c22;
               Y_7_c23 <= Y_7_c22;
               Y_8_c23 <= Y_8_c22;
               Y_9_c23 <= Y_9_c22;
               Y_10_c23 <= Y_10_c22;
               Y_11_c23 <= Y_11_c22;
               Y_12_c23 <= Y_12_c22;
               Y_13_c23 <= Y_13_c22;
               Y_14_c23 <= Y_14_c22;
               Y_15_c23 <= Y_15_c22;
               Y_16_c23 <= Y_16_c22;
               Y_17_c23 <= Y_17_c22;
               Y_18_c23 <= Y_18_c22;
               Y_19_c23 <= Y_19_c22;
               Y_20_c23 <= Y_20_c22;
               Y_21_c23 <= Y_21_c22;
               Y_22_c23 <= Y_22_c22;
            end if;
            if ce_24 = '1' then
               Y_1_c24 <= Y_1_c23;
               Y_2_c24 <= Y_2_c23;
               Y_3_c24 <= Y_3_c23;
               Y_4_c24 <= Y_4_c23;
               Y_5_c24 <= Y_5_c23;
               Y_6_c24 <= Y_6_c23;
               Y_7_c24 <= Y_7_c23;
               Y_8_c24 <= Y_8_c23;
               Y_9_c24 <= Y_9_c23;
               Y_10_c24 <= Y_10_c23;
               Y_11_c24 <= Y_11_c23;
               Y_12_c24 <= Y_12_c23;
               Y_13_c24 <= Y_13_c23;
               Y_14_c24 <= Y_14_c23;
               Y_15_c24 <= Y_15_c23;
               Y_16_c24 <= Y_16_c23;
               Y_17_c24 <= Y_17_c23;
               Y_18_c24 <= Y_18_c23;
               Y_19_c24 <= Y_19_c23;
               Y_20_c24 <= Y_20_c23;
               Y_21_c24 <= Y_21_c23;
               Y_22_c24 <= Y_22_c23;
            end if;
            if ce_25 = '1' then
               Y_1_c25 <= Y_1_c24;
               Y_2_c25 <= Y_2_c24;
               Y_3_c25 <= Y_3_c24;
               Y_4_c25 <= Y_4_c24;
               Y_5_c25 <= Y_5_c24;
               Y_6_c25 <= Y_6_c24;
               Y_7_c25 <= Y_7_c24;
               Y_8_c25 <= Y_8_c24;
               Y_9_c25 <= Y_9_c24;
               Y_10_c25 <= Y_10_c24;
               Y_11_c25 <= Y_11_c24;
               Y_12_c25 <= Y_12_c24;
               Y_13_c25 <= Y_13_c24;
               Y_14_c25 <= Y_14_c24;
               Y_15_c25 <= Y_15_c24;
               Y_16_c25 <= Y_16_c24;
               Y_17_c25 <= Y_17_c24;
               Y_18_c25 <= Y_18_c24;
               Y_19_c25 <= Y_19_c24;
               Y_20_c25 <= Y_20_c24;
               Y_21_c25 <= Y_21_c24;
               Y_22_c25 <= Y_22_c24;
            end if;
            if ce_26 = '1' then
               Y_1_c26 <= Y_1_c25;
               Y_2_c26 <= Y_2_c25;
               Y_3_c26 <= Y_3_c25;
               Y_4_c26 <= Y_4_c25;
               Y_5_c26 <= Y_5_c25;
               Y_6_c26 <= Y_6_c25;
               Y_7_c26 <= Y_7_c25;
               Y_8_c26 <= Y_8_c25;
               Y_9_c26 <= Y_9_c25;
               Y_10_c26 <= Y_10_c25;
               Y_11_c26 <= Y_11_c25;
               Y_12_c26 <= Y_12_c25;
               Y_13_c26 <= Y_13_c25;
               Y_14_c26 <= Y_14_c25;
               Y_15_c26 <= Y_15_c25;
               Y_16_c26 <= Y_16_c25;
               Y_17_c26 <= Y_17_c25;
               Y_18_c26 <= Y_18_c25;
               Y_19_c26 <= Y_19_c25;
               Y_20_c26 <= Y_20_c25;
               Y_21_c26 <= Y_21_c25;
               Y_22_c26 <= Y_22_c25;
            end if;
            if ce_27 = '1' then
               Y_1_c27 <= Y_1_c26;
               Y_2_c27 <= Y_2_c26;
               Y_3_c27 <= Y_3_c26;
               Y_4_c27 <= Y_4_c26;
               Y_5_c27 <= Y_5_c26;
               Y_6_c27 <= Y_6_c26;
               Y_7_c27 <= Y_7_c26;
               Y_8_c27 <= Y_8_c26;
               Y_9_c27 <= Y_9_c26;
               Y_10_c27 <= Y_10_c26;
               Y_11_c27 <= Y_11_c26;
               Y_12_c27 <= Y_12_c26;
               Y_13_c27 <= Y_13_c26;
               Y_14_c27 <= Y_14_c26;
               Y_15_c27 <= Y_15_c26;
               Y_16_c27 <= Y_16_c26;
               Y_17_c27 <= Y_17_c26;
               Y_18_c27 <= Y_18_c26;
               Y_19_c27 <= Y_19_c26;
               Y_20_c27 <= Y_20_c26;
               Y_21_c27 <= Y_21_c26;
               Y_22_c27 <= Y_22_c26;
            end if;
            if ce_28 = '1' then
               Y_1_c28 <= Y_1_c27;
               Y_2_c28 <= Y_2_c27;
               Y_3_c28 <= Y_3_c27;
               Y_4_c28 <= Y_4_c27;
               Y_5_c28 <= Y_5_c27;
               Y_6_c28 <= Y_6_c27;
               Y_7_c28 <= Y_7_c27;
               Y_8_c28 <= Y_8_c27;
               Y_9_c28 <= Y_9_c27;
               Y_10_c28 <= Y_10_c27;
               Y_11_c28 <= Y_11_c27;
               Y_12_c28 <= Y_12_c27;
               Y_13_c28 <= Y_13_c27;
               Y_14_c28 <= Y_14_c27;
               Y_15_c28 <= Y_15_c27;
               Y_16_c28 <= Y_16_c27;
               Y_17_c28 <= Y_17_c27;
               Y_18_c28 <= Y_18_c27;
               Y_19_c28 <= Y_19_c27;
               Y_20_c28 <= Y_20_c27;
               Y_21_c28 <= Y_21_c27;
               Y_22_c28 <= Y_22_c27;
            end if;
            if ce_29 = '1' then
               Y_1_c29 <= Y_1_c28;
               Y_2_c29 <= Y_2_c28;
               Y_3_c29 <= Y_3_c28;
               Y_4_c29 <= Y_4_c28;
               Y_5_c29 <= Y_5_c28;
               Y_6_c29 <= Y_6_c28;
               Y_7_c29 <= Y_7_c28;
               Y_8_c29 <= Y_8_c28;
               Y_9_c29 <= Y_9_c28;
               Y_10_c29 <= Y_10_c28;
               Y_11_c29 <= Y_11_c28;
               Y_12_c29 <= Y_12_c28;
               Y_13_c29 <= Y_13_c28;
               Y_14_c29 <= Y_14_c28;
               Y_15_c29 <= Y_15_c28;
               Y_16_c29 <= Y_16_c28;
               Y_17_c29 <= Y_17_c28;
               Y_18_c29 <= Y_18_c28;
               Y_19_c29 <= Y_19_c28;
               Y_20_c29 <= Y_20_c28;
               Y_21_c29 <= Y_21_c28;
               Y_22_c29 <= Y_22_c28;
            end if;
            if ce_30 = '1' then
               Y_1_c30 <= Y_1_c29;
               Y_2_c30 <= Y_2_c29;
               Y_3_c30 <= Y_3_c29;
               Y_4_c30 <= Y_4_c29;
               Y_5_c30 <= Y_5_c29;
               Y_6_c30 <= Y_6_c29;
               Y_7_c30 <= Y_7_c29;
               Y_8_c30 <= Y_8_c29;
               Y_9_c30 <= Y_9_c29;
               Y_10_c30 <= Y_10_c29;
               Y_11_c30 <= Y_11_c29;
               Y_12_c30 <= Y_12_c29;
               Y_13_c30 <= Y_13_c29;
               Y_14_c30 <= Y_14_c29;
               Y_15_c30 <= Y_15_c29;
               Y_16_c30 <= Y_16_c29;
               Y_17_c30 <= Y_17_c29;
               Y_18_c30 <= Y_18_c29;
               Y_19_c30 <= Y_19_c29;
               Y_20_c30 <= Y_20_c29;
               Y_21_c30 <= Y_21_c29;
               Y_22_c30 <= Y_22_c29;
            end if;
            if ce_31 = '1' then
               Y_1_c31 <= Y_1_c30;
               Y_2_c31 <= Y_2_c30;
               Y_3_c31 <= Y_3_c30;
               Y_4_c31 <= Y_4_c30;
               Y_5_c31 <= Y_5_c30;
               Y_6_c31 <= Y_6_c30;
               Y_7_c31 <= Y_7_c30;
               Y_8_c31 <= Y_8_c30;
               Y_9_c31 <= Y_9_c30;
               Y_10_c31 <= Y_10_c30;
               Y_11_c31 <= Y_11_c30;
               Y_12_c31 <= Y_12_c30;
               Y_13_c31 <= Y_13_c30;
               Y_14_c31 <= Y_14_c30;
               Y_15_c31 <= Y_15_c30;
               Y_16_c31 <= Y_16_c30;
               Y_17_c31 <= Y_17_c30;
               Y_18_c31 <= Y_18_c30;
               Y_19_c31 <= Y_19_c30;
               Y_20_c31 <= Y_20_c30;
               Y_21_c31 <= Y_21_c30;
               Y_22_c31 <= Y_22_c30;
            end if;
            if ce_32 = '1' then
               Y_1_c32 <= Y_1_c31;
               Y_2_c32 <= Y_2_c31;
               Y_3_c32 <= Y_3_c31;
               Y_4_c32 <= Y_4_c31;
               Y_5_c32 <= Y_5_c31;
               Y_6_c32 <= Y_6_c31;
               Y_7_c32 <= Y_7_c31;
               Y_8_c32 <= Y_8_c31;
               Y_9_c32 <= Y_9_c31;
               Y_10_c32 <= Y_10_c31;
               Y_11_c32 <= Y_11_c31;
               Y_12_c32 <= Y_12_c31;
               Y_13_c32 <= Y_13_c31;
               Y_14_c32 <= Y_14_c31;
               Y_15_c32 <= Y_15_c31;
               Y_16_c32 <= Y_16_c31;
               Y_17_c32 <= Y_17_c31;
               Y_18_c32 <= Y_18_c31;
               Y_19_c32 <= Y_19_c31;
               Y_20_c32 <= Y_20_c31;
               Y_21_c32 <= Y_21_c31;
               Y_22_c32 <= Y_22_c31;
            end if;
            if ce_33 = '1' then
               Y_1_c33 <= Y_1_c32;
               Y_2_c33 <= Y_2_c32;
               Y_3_c33 <= Y_3_c32;
               Y_4_c33 <= Y_4_c32;
               Y_5_c33 <= Y_5_c32;
               Y_6_c33 <= Y_6_c32;
               Y_7_c33 <= Y_7_c32;
               Y_8_c33 <= Y_8_c32;
               Y_9_c33 <= Y_9_c32;
               Y_10_c33 <= Y_10_c32;
               Y_11_c33 <= Y_11_c32;
               Y_12_c33 <= Y_12_c32;
               Y_13_c33 <= Y_13_c32;
               Y_14_c33 <= Y_14_c32;
               Y_15_c33 <= Y_15_c32;
               Y_16_c33 <= Y_16_c32;
               Y_17_c33 <= Y_17_c32;
               Y_18_c33 <= Y_18_c32;
               Y_19_c33 <= Y_19_c32;
               Y_20_c33 <= Y_20_c32;
               Y_21_c33 <= Y_21_c32;
               Y_22_c33 <= Y_22_c32;
            end if;
            if ce_34 = '1' then
               X_1_c34 <= X_1_c33;
               Y_1_c34 <= Y_1_c33;
               X_2_c34 <= X_2_c33;
               Y_2_c34 <= Y_2_c33;
               X_3_c34 <= X_3_c33;
               Y_3_c34 <= Y_3_c33;
               X_4_c34 <= X_4_c33;
               Y_4_c34 <= Y_4_c33;
               X_5_c34 <= X_5_c33;
               Y_5_c34 <= Y_5_c33;
               X_6_c34 <= X_6_c33;
               Y_6_c34 <= Y_6_c33;
               X_7_c34 <= X_7_c33;
               Y_7_c34 <= Y_7_c33;
               X_8_c34 <= X_8_c33;
               Y_8_c34 <= Y_8_c33;
               X_9_c34 <= X_9_c33;
               Y_9_c34 <= Y_9_c33;
               X_10_c34 <= X_10_c33;
               Y_10_c34 <= Y_10_c33;
               X_11_c34 <= X_11_c33;
               Y_11_c34 <= Y_11_c33;
               X_12_c34 <= X_12_c33;
               Y_12_c34 <= Y_12_c33;
               X_13_c34 <= X_13_c33;
               Y_13_c34 <= Y_13_c33;
               X_14_c34 <= X_14_c33;
               Y_14_c34 <= Y_14_c33;
               X_15_c34 <= X_15_c33;
               Y_15_c34 <= Y_15_c33;
               X_16_c34 <= X_16_c33;
               Y_16_c34 <= Y_16_c33;
               X_17_c34 <= X_17_c33;
               Y_17_c34 <= Y_17_c33;
               X_18_c34 <= X_18_c33;
               Y_18_c34 <= Y_18_c33;
               X_19_c34 <= X_19_c33;
               Y_19_c34 <= Y_19_c33;
               X_20_c34 <= X_20_c33;
               Y_20_c34 <= Y_20_c33;
               X_21_c34 <= X_21_c33;
               Y_21_c34 <= Y_21_c33;
               X_22_c34 <= X_22_c33;
               Y_22_c34 <= Y_22_c33;
            end if;
            if ce_35 = '1' then
               Cin_1_c35 <= Cin_1_c34;
               X_1_c35 <= X_1_c34;
               Y_1_c35 <= Y_1_c34;
               X_2_c35 <= X_2_c34;
               Y_2_c35 <= Y_2_c34;
               X_3_c35 <= X_3_c34;
               Y_3_c35 <= Y_3_c34;
               X_4_c35 <= X_4_c34;
               Y_4_c35 <= Y_4_c34;
               X_5_c35 <= X_5_c34;
               Y_5_c35 <= Y_5_c34;
               X_6_c35 <= X_6_c34;
               Y_6_c35 <= Y_6_c34;
               X_7_c35 <= X_7_c34;
               Y_7_c35 <= Y_7_c34;
               X_8_c35 <= X_8_c34;
               Y_8_c35 <= Y_8_c34;
               X_9_c35 <= X_9_c34;
               Y_9_c35 <= Y_9_c34;
               X_10_c35 <= X_10_c34;
               Y_10_c35 <= Y_10_c34;
               X_11_c35 <= X_11_c34;
               Y_11_c35 <= Y_11_c34;
               X_12_c35 <= X_12_c34;
               Y_12_c35 <= Y_12_c34;
               X_13_c35 <= X_13_c34;
               Y_13_c35 <= Y_13_c34;
               X_14_c35 <= X_14_c34;
               Y_14_c35 <= Y_14_c34;
               X_15_c35 <= X_15_c34;
               Y_15_c35 <= Y_15_c34;
               X_16_c35 <= X_16_c34;
               Y_16_c35 <= Y_16_c34;
               X_17_c35 <= X_17_c34;
               Y_17_c35 <= Y_17_c34;
               X_18_c35 <= X_18_c34;
               Y_18_c35 <= Y_18_c34;
               X_19_c35 <= X_19_c34;
               Y_19_c35 <= Y_19_c34;
               X_20_c35 <= X_20_c34;
               Y_20_c35 <= Y_20_c34;
               X_21_c35 <= X_21_c34;
               Y_21_c35 <= Y_21_c34;
               X_22_c35 <= X_22_c34;
               Y_22_c35 <= Y_22_c34;
            end if;
            if ce_36 = '1' then
               R_1_c36 <= R_1_c35;
               Cin_2_c36 <= Cin_2_c35;
               X_2_c36 <= X_2_c35;
               Y_2_c36 <= Y_2_c35;
               X_3_c36 <= X_3_c35;
               Y_3_c36 <= Y_3_c35;
               X_4_c36 <= X_4_c35;
               Y_4_c36 <= Y_4_c35;
               X_5_c36 <= X_5_c35;
               Y_5_c36 <= Y_5_c35;
               X_6_c36 <= X_6_c35;
               Y_6_c36 <= Y_6_c35;
               X_7_c36 <= X_7_c35;
               Y_7_c36 <= Y_7_c35;
               X_8_c36 <= X_8_c35;
               Y_8_c36 <= Y_8_c35;
               X_9_c36 <= X_9_c35;
               Y_9_c36 <= Y_9_c35;
               X_10_c36 <= X_10_c35;
               Y_10_c36 <= Y_10_c35;
               X_11_c36 <= X_11_c35;
               Y_11_c36 <= Y_11_c35;
               X_12_c36 <= X_12_c35;
               Y_12_c36 <= Y_12_c35;
               X_13_c36 <= X_13_c35;
               Y_13_c36 <= Y_13_c35;
               X_14_c36 <= X_14_c35;
               Y_14_c36 <= Y_14_c35;
               X_15_c36 <= X_15_c35;
               Y_15_c36 <= Y_15_c35;
               X_16_c36 <= X_16_c35;
               Y_16_c36 <= Y_16_c35;
               X_17_c36 <= X_17_c35;
               Y_17_c36 <= Y_17_c35;
               X_18_c36 <= X_18_c35;
               Y_18_c36 <= Y_18_c35;
               X_19_c36 <= X_19_c35;
               Y_19_c36 <= Y_19_c35;
               X_20_c36 <= X_20_c35;
               Y_20_c36 <= Y_20_c35;
               X_21_c36 <= X_21_c35;
               Y_21_c36 <= Y_21_c35;
               X_22_c36 <= X_22_c35;
               Y_22_c36 <= Y_22_c35;
            end if;
            if ce_37 = '1' then
               R_1_c37 <= R_1_c36;
               R_2_c37 <= R_2_c36;
               Cin_3_c37 <= Cin_3_c36;
               X_3_c37 <= X_3_c36;
               Y_3_c37 <= Y_3_c36;
               X_4_c37 <= X_4_c36;
               Y_4_c37 <= Y_4_c36;
               X_5_c37 <= X_5_c36;
               Y_5_c37 <= Y_5_c36;
               X_6_c37 <= X_6_c36;
               Y_6_c37 <= Y_6_c36;
               X_7_c37 <= X_7_c36;
               Y_7_c37 <= Y_7_c36;
               X_8_c37 <= X_8_c36;
               Y_8_c37 <= Y_8_c36;
               X_9_c37 <= X_9_c36;
               Y_9_c37 <= Y_9_c36;
               X_10_c37 <= X_10_c36;
               Y_10_c37 <= Y_10_c36;
               X_11_c37 <= X_11_c36;
               Y_11_c37 <= Y_11_c36;
               X_12_c37 <= X_12_c36;
               Y_12_c37 <= Y_12_c36;
               X_13_c37 <= X_13_c36;
               Y_13_c37 <= Y_13_c36;
               X_14_c37 <= X_14_c36;
               Y_14_c37 <= Y_14_c36;
               X_15_c37 <= X_15_c36;
               Y_15_c37 <= Y_15_c36;
               X_16_c37 <= X_16_c36;
               Y_16_c37 <= Y_16_c36;
               X_17_c37 <= X_17_c36;
               Y_17_c37 <= Y_17_c36;
               X_18_c37 <= X_18_c36;
               Y_18_c37 <= Y_18_c36;
               X_19_c37 <= X_19_c36;
               Y_19_c37 <= Y_19_c36;
               X_20_c37 <= X_20_c36;
               Y_20_c37 <= Y_20_c36;
               X_21_c37 <= X_21_c36;
               Y_21_c37 <= Y_21_c36;
               X_22_c37 <= X_22_c36;
               Y_22_c37 <= Y_22_c36;
            end if;
            if ce_38 = '1' then
               R_1_c38 <= R_1_c37;
               R_2_c38 <= R_2_c37;
               R_3_c38 <= R_3_c37;
               Cin_4_c38 <= Cin_4_c37;
               X_4_c38 <= X_4_c37;
               Y_4_c38 <= Y_4_c37;
               X_5_c38 <= X_5_c37;
               Y_5_c38 <= Y_5_c37;
               X_6_c38 <= X_6_c37;
               Y_6_c38 <= Y_6_c37;
               X_7_c38 <= X_7_c37;
               Y_7_c38 <= Y_7_c37;
               X_8_c38 <= X_8_c37;
               Y_8_c38 <= Y_8_c37;
               X_9_c38 <= X_9_c37;
               Y_9_c38 <= Y_9_c37;
               X_10_c38 <= X_10_c37;
               Y_10_c38 <= Y_10_c37;
               X_11_c38 <= X_11_c37;
               Y_11_c38 <= Y_11_c37;
               X_12_c38 <= X_12_c37;
               Y_12_c38 <= Y_12_c37;
               X_13_c38 <= X_13_c37;
               Y_13_c38 <= Y_13_c37;
               X_14_c38 <= X_14_c37;
               Y_14_c38 <= Y_14_c37;
               X_15_c38 <= X_15_c37;
               Y_15_c38 <= Y_15_c37;
               X_16_c38 <= X_16_c37;
               Y_16_c38 <= Y_16_c37;
               X_17_c38 <= X_17_c37;
               Y_17_c38 <= Y_17_c37;
               X_18_c38 <= X_18_c37;
               Y_18_c38 <= Y_18_c37;
               X_19_c38 <= X_19_c37;
               Y_19_c38 <= Y_19_c37;
               X_20_c38 <= X_20_c37;
               Y_20_c38 <= Y_20_c37;
               X_21_c38 <= X_21_c37;
               Y_21_c38 <= Y_21_c37;
               X_22_c38 <= X_22_c37;
               Y_22_c38 <= Y_22_c37;
            end if;
            if ce_39 = '1' then
               R_1_c39 <= R_1_c38;
               R_2_c39 <= R_2_c38;
               R_3_c39 <= R_3_c38;
               R_4_c39 <= R_4_c38;
               Cin_5_c39 <= Cin_5_c38;
               X_5_c39 <= X_5_c38;
               Y_5_c39 <= Y_5_c38;
               X_6_c39 <= X_6_c38;
               Y_6_c39 <= Y_6_c38;
               X_7_c39 <= X_7_c38;
               Y_7_c39 <= Y_7_c38;
               X_8_c39 <= X_8_c38;
               Y_8_c39 <= Y_8_c38;
               X_9_c39 <= X_9_c38;
               Y_9_c39 <= Y_9_c38;
               X_10_c39 <= X_10_c38;
               Y_10_c39 <= Y_10_c38;
               X_11_c39 <= X_11_c38;
               Y_11_c39 <= Y_11_c38;
               X_12_c39 <= X_12_c38;
               Y_12_c39 <= Y_12_c38;
               X_13_c39 <= X_13_c38;
               Y_13_c39 <= Y_13_c38;
               X_14_c39 <= X_14_c38;
               Y_14_c39 <= Y_14_c38;
               X_15_c39 <= X_15_c38;
               Y_15_c39 <= Y_15_c38;
               X_16_c39 <= X_16_c38;
               Y_16_c39 <= Y_16_c38;
               X_17_c39 <= X_17_c38;
               Y_17_c39 <= Y_17_c38;
               X_18_c39 <= X_18_c38;
               Y_18_c39 <= Y_18_c38;
               X_19_c39 <= X_19_c38;
               Y_19_c39 <= Y_19_c38;
               X_20_c39 <= X_20_c38;
               Y_20_c39 <= Y_20_c38;
               X_21_c39 <= X_21_c38;
               Y_21_c39 <= Y_21_c38;
               X_22_c39 <= X_22_c38;
               Y_22_c39 <= Y_22_c38;
            end if;
            if ce_40 = '1' then
               R_1_c40 <= R_1_c39;
               R_2_c40 <= R_2_c39;
               R_3_c40 <= R_3_c39;
               R_4_c40 <= R_4_c39;
               R_5_c40 <= R_5_c39;
               Cin_6_c40 <= Cin_6_c39;
               X_6_c40 <= X_6_c39;
               Y_6_c40 <= Y_6_c39;
               X_7_c40 <= X_7_c39;
               Y_7_c40 <= Y_7_c39;
               X_8_c40 <= X_8_c39;
               Y_8_c40 <= Y_8_c39;
               X_9_c40 <= X_9_c39;
               Y_9_c40 <= Y_9_c39;
               X_10_c40 <= X_10_c39;
               Y_10_c40 <= Y_10_c39;
               X_11_c40 <= X_11_c39;
               Y_11_c40 <= Y_11_c39;
               X_12_c40 <= X_12_c39;
               Y_12_c40 <= Y_12_c39;
               X_13_c40 <= X_13_c39;
               Y_13_c40 <= Y_13_c39;
               X_14_c40 <= X_14_c39;
               Y_14_c40 <= Y_14_c39;
               X_15_c40 <= X_15_c39;
               Y_15_c40 <= Y_15_c39;
               X_16_c40 <= X_16_c39;
               Y_16_c40 <= Y_16_c39;
               X_17_c40 <= X_17_c39;
               Y_17_c40 <= Y_17_c39;
               X_18_c40 <= X_18_c39;
               Y_18_c40 <= Y_18_c39;
               X_19_c40 <= X_19_c39;
               Y_19_c40 <= Y_19_c39;
               X_20_c40 <= X_20_c39;
               Y_20_c40 <= Y_20_c39;
               X_21_c40 <= X_21_c39;
               Y_21_c40 <= Y_21_c39;
               X_22_c40 <= X_22_c39;
               Y_22_c40 <= Y_22_c39;
            end if;
            if ce_41 = '1' then
               R_1_c41 <= R_1_c40;
               R_2_c41 <= R_2_c40;
               R_3_c41 <= R_3_c40;
               R_4_c41 <= R_4_c40;
               R_5_c41 <= R_5_c40;
               R_6_c41 <= R_6_c40;
               Cin_7_c41 <= Cin_7_c40;
               X_7_c41 <= X_7_c40;
               Y_7_c41 <= Y_7_c40;
               X_8_c41 <= X_8_c40;
               Y_8_c41 <= Y_8_c40;
               X_9_c41 <= X_9_c40;
               Y_9_c41 <= Y_9_c40;
               X_10_c41 <= X_10_c40;
               Y_10_c41 <= Y_10_c40;
               X_11_c41 <= X_11_c40;
               Y_11_c41 <= Y_11_c40;
               X_12_c41 <= X_12_c40;
               Y_12_c41 <= Y_12_c40;
               X_13_c41 <= X_13_c40;
               Y_13_c41 <= Y_13_c40;
               X_14_c41 <= X_14_c40;
               Y_14_c41 <= Y_14_c40;
               X_15_c41 <= X_15_c40;
               Y_15_c41 <= Y_15_c40;
               X_16_c41 <= X_16_c40;
               Y_16_c41 <= Y_16_c40;
               X_17_c41 <= X_17_c40;
               Y_17_c41 <= Y_17_c40;
               X_18_c41 <= X_18_c40;
               Y_18_c41 <= Y_18_c40;
               X_19_c41 <= X_19_c40;
               Y_19_c41 <= Y_19_c40;
               X_20_c41 <= X_20_c40;
               Y_20_c41 <= Y_20_c40;
               X_21_c41 <= X_21_c40;
               Y_21_c41 <= Y_21_c40;
               X_22_c41 <= X_22_c40;
               Y_22_c41 <= Y_22_c40;
            end if;
            if ce_42 = '1' then
               R_1_c42 <= R_1_c41;
               R_2_c42 <= R_2_c41;
               R_3_c42 <= R_3_c41;
               R_4_c42 <= R_4_c41;
               R_5_c42 <= R_5_c41;
               R_6_c42 <= R_6_c41;
               R_7_c42 <= R_7_c41;
               Cin_8_c42 <= Cin_8_c41;
               X_8_c42 <= X_8_c41;
               Y_8_c42 <= Y_8_c41;
               X_9_c42 <= X_9_c41;
               Y_9_c42 <= Y_9_c41;
               X_10_c42 <= X_10_c41;
               Y_10_c42 <= Y_10_c41;
               X_11_c42 <= X_11_c41;
               Y_11_c42 <= Y_11_c41;
               X_12_c42 <= X_12_c41;
               Y_12_c42 <= Y_12_c41;
               X_13_c42 <= X_13_c41;
               Y_13_c42 <= Y_13_c41;
               X_14_c42 <= X_14_c41;
               Y_14_c42 <= Y_14_c41;
               X_15_c42 <= X_15_c41;
               Y_15_c42 <= Y_15_c41;
               X_16_c42 <= X_16_c41;
               Y_16_c42 <= Y_16_c41;
               X_17_c42 <= X_17_c41;
               Y_17_c42 <= Y_17_c41;
               X_18_c42 <= X_18_c41;
               Y_18_c42 <= Y_18_c41;
               X_19_c42 <= X_19_c41;
               Y_19_c42 <= Y_19_c41;
               X_20_c42 <= X_20_c41;
               Y_20_c42 <= Y_20_c41;
               X_21_c42 <= X_21_c41;
               Y_21_c42 <= Y_21_c41;
               X_22_c42 <= X_22_c41;
               Y_22_c42 <= Y_22_c41;
            end if;
            if ce_43 = '1' then
               R_1_c43 <= R_1_c42;
               R_2_c43 <= R_2_c42;
               R_3_c43 <= R_3_c42;
               R_4_c43 <= R_4_c42;
               R_5_c43 <= R_5_c42;
               R_6_c43 <= R_6_c42;
               R_7_c43 <= R_7_c42;
               R_8_c43 <= R_8_c42;
               Cin_9_c43 <= Cin_9_c42;
               X_9_c43 <= X_9_c42;
               Y_9_c43 <= Y_9_c42;
               X_10_c43 <= X_10_c42;
               Y_10_c43 <= Y_10_c42;
               X_11_c43 <= X_11_c42;
               Y_11_c43 <= Y_11_c42;
               X_12_c43 <= X_12_c42;
               Y_12_c43 <= Y_12_c42;
               X_13_c43 <= X_13_c42;
               Y_13_c43 <= Y_13_c42;
               X_14_c43 <= X_14_c42;
               Y_14_c43 <= Y_14_c42;
               X_15_c43 <= X_15_c42;
               Y_15_c43 <= Y_15_c42;
               X_16_c43 <= X_16_c42;
               Y_16_c43 <= Y_16_c42;
               X_17_c43 <= X_17_c42;
               Y_17_c43 <= Y_17_c42;
               X_18_c43 <= X_18_c42;
               Y_18_c43 <= Y_18_c42;
               X_19_c43 <= X_19_c42;
               Y_19_c43 <= Y_19_c42;
               X_20_c43 <= X_20_c42;
               Y_20_c43 <= Y_20_c42;
               X_21_c43 <= X_21_c42;
               Y_21_c43 <= Y_21_c42;
               X_22_c43 <= X_22_c42;
               Y_22_c43 <= Y_22_c42;
            end if;
            if ce_44 = '1' then
               R_1_c44 <= R_1_c43;
               R_2_c44 <= R_2_c43;
               R_3_c44 <= R_3_c43;
               R_4_c44 <= R_4_c43;
               R_5_c44 <= R_5_c43;
               R_6_c44 <= R_6_c43;
               R_7_c44 <= R_7_c43;
               R_8_c44 <= R_8_c43;
               R_9_c44 <= R_9_c43;
               Cin_10_c44 <= Cin_10_c43;
               X_10_c44 <= X_10_c43;
               Y_10_c44 <= Y_10_c43;
               X_11_c44 <= X_11_c43;
               Y_11_c44 <= Y_11_c43;
               X_12_c44 <= X_12_c43;
               Y_12_c44 <= Y_12_c43;
               X_13_c44 <= X_13_c43;
               Y_13_c44 <= Y_13_c43;
               X_14_c44 <= X_14_c43;
               Y_14_c44 <= Y_14_c43;
               X_15_c44 <= X_15_c43;
               Y_15_c44 <= Y_15_c43;
               X_16_c44 <= X_16_c43;
               Y_16_c44 <= Y_16_c43;
               X_17_c44 <= X_17_c43;
               Y_17_c44 <= Y_17_c43;
               X_18_c44 <= X_18_c43;
               Y_18_c44 <= Y_18_c43;
               X_19_c44 <= X_19_c43;
               Y_19_c44 <= Y_19_c43;
               X_20_c44 <= X_20_c43;
               Y_20_c44 <= Y_20_c43;
               X_21_c44 <= X_21_c43;
               Y_21_c44 <= Y_21_c43;
               X_22_c44 <= X_22_c43;
               Y_22_c44 <= Y_22_c43;
            end if;
            if ce_45 = '1' then
               R_1_c45 <= R_1_c44;
               R_2_c45 <= R_2_c44;
               R_3_c45 <= R_3_c44;
               R_4_c45 <= R_4_c44;
               R_5_c45 <= R_5_c44;
               R_6_c45 <= R_6_c44;
               R_7_c45 <= R_7_c44;
               R_8_c45 <= R_8_c44;
               R_9_c45 <= R_9_c44;
               R_10_c45 <= R_10_c44;
               Cin_11_c45 <= Cin_11_c44;
               X_11_c45 <= X_11_c44;
               Y_11_c45 <= Y_11_c44;
               X_12_c45 <= X_12_c44;
               Y_12_c45 <= Y_12_c44;
               X_13_c45 <= X_13_c44;
               Y_13_c45 <= Y_13_c44;
               X_14_c45 <= X_14_c44;
               Y_14_c45 <= Y_14_c44;
               X_15_c45 <= X_15_c44;
               Y_15_c45 <= Y_15_c44;
               X_16_c45 <= X_16_c44;
               Y_16_c45 <= Y_16_c44;
               X_17_c45 <= X_17_c44;
               Y_17_c45 <= Y_17_c44;
               X_18_c45 <= X_18_c44;
               Y_18_c45 <= Y_18_c44;
               X_19_c45 <= X_19_c44;
               Y_19_c45 <= Y_19_c44;
               X_20_c45 <= X_20_c44;
               Y_20_c45 <= Y_20_c44;
               X_21_c45 <= X_21_c44;
               Y_21_c45 <= Y_21_c44;
               X_22_c45 <= X_22_c44;
               Y_22_c45 <= Y_22_c44;
            end if;
            if ce_46 = '1' then
               R_1_c46 <= R_1_c45;
               R_2_c46 <= R_2_c45;
               R_3_c46 <= R_3_c45;
               R_4_c46 <= R_4_c45;
               R_5_c46 <= R_5_c45;
               R_6_c46 <= R_6_c45;
               R_7_c46 <= R_7_c45;
               R_8_c46 <= R_8_c45;
               R_9_c46 <= R_9_c45;
               R_10_c46 <= R_10_c45;
               R_11_c46 <= R_11_c45;
               Cin_12_c46 <= Cin_12_c45;
               X_12_c46 <= X_12_c45;
               Y_12_c46 <= Y_12_c45;
               X_13_c46 <= X_13_c45;
               Y_13_c46 <= Y_13_c45;
               X_14_c46 <= X_14_c45;
               Y_14_c46 <= Y_14_c45;
               X_15_c46 <= X_15_c45;
               Y_15_c46 <= Y_15_c45;
               X_16_c46 <= X_16_c45;
               Y_16_c46 <= Y_16_c45;
               X_17_c46 <= X_17_c45;
               Y_17_c46 <= Y_17_c45;
               X_18_c46 <= X_18_c45;
               Y_18_c46 <= Y_18_c45;
               X_19_c46 <= X_19_c45;
               Y_19_c46 <= Y_19_c45;
               X_20_c46 <= X_20_c45;
               Y_20_c46 <= Y_20_c45;
               X_21_c46 <= X_21_c45;
               Y_21_c46 <= Y_21_c45;
               X_22_c46 <= X_22_c45;
               Y_22_c46 <= Y_22_c45;
            end if;
            if ce_47 = '1' then
               R_1_c47 <= R_1_c46;
               R_2_c47 <= R_2_c46;
               R_3_c47 <= R_3_c46;
               R_4_c47 <= R_4_c46;
               R_5_c47 <= R_5_c46;
               R_6_c47 <= R_6_c46;
               R_7_c47 <= R_7_c46;
               R_8_c47 <= R_8_c46;
               R_9_c47 <= R_9_c46;
               R_10_c47 <= R_10_c46;
               R_11_c47 <= R_11_c46;
               R_12_c47 <= R_12_c46;
               Cin_13_c47 <= Cin_13_c46;
               X_13_c47 <= X_13_c46;
               Y_13_c47 <= Y_13_c46;
               X_14_c47 <= X_14_c46;
               Y_14_c47 <= Y_14_c46;
               X_15_c47 <= X_15_c46;
               Y_15_c47 <= Y_15_c46;
               X_16_c47 <= X_16_c46;
               Y_16_c47 <= Y_16_c46;
               X_17_c47 <= X_17_c46;
               Y_17_c47 <= Y_17_c46;
               X_18_c47 <= X_18_c46;
               Y_18_c47 <= Y_18_c46;
               X_19_c47 <= X_19_c46;
               Y_19_c47 <= Y_19_c46;
               X_20_c47 <= X_20_c46;
               Y_20_c47 <= Y_20_c46;
               X_21_c47 <= X_21_c46;
               Y_21_c47 <= Y_21_c46;
               X_22_c47 <= X_22_c46;
               Y_22_c47 <= Y_22_c46;
            end if;
            if ce_48 = '1' then
               R_1_c48 <= R_1_c47;
               R_2_c48 <= R_2_c47;
               R_3_c48 <= R_3_c47;
               R_4_c48 <= R_4_c47;
               R_5_c48 <= R_5_c47;
               R_6_c48 <= R_6_c47;
               R_7_c48 <= R_7_c47;
               R_8_c48 <= R_8_c47;
               R_9_c48 <= R_9_c47;
               R_10_c48 <= R_10_c47;
               R_11_c48 <= R_11_c47;
               R_12_c48 <= R_12_c47;
               R_13_c48 <= R_13_c47;
               Cin_14_c48 <= Cin_14_c47;
               X_14_c48 <= X_14_c47;
               Y_14_c48 <= Y_14_c47;
               X_15_c48 <= X_15_c47;
               Y_15_c48 <= Y_15_c47;
               X_16_c48 <= X_16_c47;
               Y_16_c48 <= Y_16_c47;
               X_17_c48 <= X_17_c47;
               Y_17_c48 <= Y_17_c47;
               X_18_c48 <= X_18_c47;
               Y_18_c48 <= Y_18_c47;
               X_19_c48 <= X_19_c47;
               Y_19_c48 <= Y_19_c47;
               X_20_c48 <= X_20_c47;
               Y_20_c48 <= Y_20_c47;
               X_21_c48 <= X_21_c47;
               Y_21_c48 <= Y_21_c47;
               X_22_c48 <= X_22_c47;
               Y_22_c48 <= Y_22_c47;
            end if;
            if ce_49 = '1' then
               R_1_c49 <= R_1_c48;
               R_2_c49 <= R_2_c48;
               R_3_c49 <= R_3_c48;
               R_4_c49 <= R_4_c48;
               R_5_c49 <= R_5_c48;
               R_6_c49 <= R_6_c48;
               R_7_c49 <= R_7_c48;
               R_8_c49 <= R_8_c48;
               R_9_c49 <= R_9_c48;
               R_10_c49 <= R_10_c48;
               R_11_c49 <= R_11_c48;
               R_12_c49 <= R_12_c48;
               R_13_c49 <= R_13_c48;
               R_14_c49 <= R_14_c48;
               Cin_15_c49 <= Cin_15_c48;
               X_15_c49 <= X_15_c48;
               Y_15_c49 <= Y_15_c48;
               X_16_c49 <= X_16_c48;
               Y_16_c49 <= Y_16_c48;
               X_17_c49 <= X_17_c48;
               Y_17_c49 <= Y_17_c48;
               X_18_c49 <= X_18_c48;
               Y_18_c49 <= Y_18_c48;
               X_19_c49 <= X_19_c48;
               Y_19_c49 <= Y_19_c48;
               X_20_c49 <= X_20_c48;
               Y_20_c49 <= Y_20_c48;
               X_21_c49 <= X_21_c48;
               Y_21_c49 <= Y_21_c48;
               X_22_c49 <= X_22_c48;
               Y_22_c49 <= Y_22_c48;
            end if;
            if ce_50 = '1' then
               R_1_c50 <= R_1_c49;
               R_2_c50 <= R_2_c49;
               R_3_c50 <= R_3_c49;
               R_4_c50 <= R_4_c49;
               R_5_c50 <= R_5_c49;
               R_6_c50 <= R_6_c49;
               R_7_c50 <= R_7_c49;
               R_8_c50 <= R_8_c49;
               R_9_c50 <= R_9_c49;
               R_10_c50 <= R_10_c49;
               R_11_c50 <= R_11_c49;
               R_12_c50 <= R_12_c49;
               R_13_c50 <= R_13_c49;
               R_14_c50 <= R_14_c49;
               R_15_c50 <= R_15_c49;
               Cin_16_c50 <= Cin_16_c49;
               X_16_c50 <= X_16_c49;
               Y_16_c50 <= Y_16_c49;
               X_17_c50 <= X_17_c49;
               Y_17_c50 <= Y_17_c49;
               X_18_c50 <= X_18_c49;
               Y_18_c50 <= Y_18_c49;
               X_19_c50 <= X_19_c49;
               Y_19_c50 <= Y_19_c49;
               X_20_c50 <= X_20_c49;
               Y_20_c50 <= Y_20_c49;
               X_21_c50 <= X_21_c49;
               Y_21_c50 <= Y_21_c49;
               X_22_c50 <= X_22_c49;
               Y_22_c50 <= Y_22_c49;
            end if;
            if ce_51 = '1' then
               R_1_c51 <= R_1_c50;
               R_2_c51 <= R_2_c50;
               R_3_c51 <= R_3_c50;
               R_4_c51 <= R_4_c50;
               R_5_c51 <= R_5_c50;
               R_6_c51 <= R_6_c50;
               R_7_c51 <= R_7_c50;
               R_8_c51 <= R_8_c50;
               R_9_c51 <= R_9_c50;
               R_10_c51 <= R_10_c50;
               R_11_c51 <= R_11_c50;
               R_12_c51 <= R_12_c50;
               R_13_c51 <= R_13_c50;
               R_14_c51 <= R_14_c50;
               R_15_c51 <= R_15_c50;
               R_16_c51 <= R_16_c50;
               Cin_17_c51 <= Cin_17_c50;
               X_17_c51 <= X_17_c50;
               Y_17_c51 <= Y_17_c50;
               X_18_c51 <= X_18_c50;
               Y_18_c51 <= Y_18_c50;
               X_19_c51 <= X_19_c50;
               Y_19_c51 <= Y_19_c50;
               X_20_c51 <= X_20_c50;
               Y_20_c51 <= Y_20_c50;
               X_21_c51 <= X_21_c50;
               Y_21_c51 <= Y_21_c50;
               X_22_c51 <= X_22_c50;
               Y_22_c51 <= Y_22_c50;
            end if;
            if ce_52 = '1' then
               R_1_c52 <= R_1_c51;
               R_2_c52 <= R_2_c51;
               R_3_c52 <= R_3_c51;
               R_4_c52 <= R_4_c51;
               R_5_c52 <= R_5_c51;
               R_6_c52 <= R_6_c51;
               R_7_c52 <= R_7_c51;
               R_8_c52 <= R_8_c51;
               R_9_c52 <= R_9_c51;
               R_10_c52 <= R_10_c51;
               R_11_c52 <= R_11_c51;
               R_12_c52 <= R_12_c51;
               R_13_c52 <= R_13_c51;
               R_14_c52 <= R_14_c51;
               R_15_c52 <= R_15_c51;
               R_16_c52 <= R_16_c51;
               R_17_c52 <= R_17_c51;
               Cin_18_c52 <= Cin_18_c51;
               X_18_c52 <= X_18_c51;
               Y_18_c52 <= Y_18_c51;
               X_19_c52 <= X_19_c51;
               Y_19_c52 <= Y_19_c51;
               X_20_c52 <= X_20_c51;
               Y_20_c52 <= Y_20_c51;
               X_21_c52 <= X_21_c51;
               Y_21_c52 <= Y_21_c51;
               X_22_c52 <= X_22_c51;
               Y_22_c52 <= Y_22_c51;
            end if;
            if ce_53 = '1' then
               R_1_c53 <= R_1_c52;
               R_2_c53 <= R_2_c52;
               R_3_c53 <= R_3_c52;
               R_4_c53 <= R_4_c52;
               R_5_c53 <= R_5_c52;
               R_6_c53 <= R_6_c52;
               R_7_c53 <= R_7_c52;
               R_8_c53 <= R_8_c52;
               R_9_c53 <= R_9_c52;
               R_10_c53 <= R_10_c52;
               R_11_c53 <= R_11_c52;
               R_12_c53 <= R_12_c52;
               R_13_c53 <= R_13_c52;
               R_14_c53 <= R_14_c52;
               R_15_c53 <= R_15_c52;
               R_16_c53 <= R_16_c52;
               R_17_c53 <= R_17_c52;
               R_18_c53 <= R_18_c52;
               Cin_19_c53 <= Cin_19_c52;
               X_19_c53 <= X_19_c52;
               Y_19_c53 <= Y_19_c52;
               X_20_c53 <= X_20_c52;
               Y_20_c53 <= Y_20_c52;
               X_21_c53 <= X_21_c52;
               Y_21_c53 <= Y_21_c52;
               X_22_c53 <= X_22_c52;
               Y_22_c53 <= Y_22_c52;
            end if;
            if ce_54 = '1' then
               R_1_c54 <= R_1_c53;
               R_2_c54 <= R_2_c53;
               R_3_c54 <= R_3_c53;
               R_4_c54 <= R_4_c53;
               R_5_c54 <= R_5_c53;
               R_6_c54 <= R_6_c53;
               R_7_c54 <= R_7_c53;
               R_8_c54 <= R_8_c53;
               R_9_c54 <= R_9_c53;
               R_10_c54 <= R_10_c53;
               R_11_c54 <= R_11_c53;
               R_12_c54 <= R_12_c53;
               R_13_c54 <= R_13_c53;
               R_14_c54 <= R_14_c53;
               R_15_c54 <= R_15_c53;
               R_16_c54 <= R_16_c53;
               R_17_c54 <= R_17_c53;
               R_18_c54 <= R_18_c53;
               R_19_c54 <= R_19_c53;
               Cin_20_c54 <= Cin_20_c53;
               X_20_c54 <= X_20_c53;
               Y_20_c54 <= Y_20_c53;
               X_21_c54 <= X_21_c53;
               Y_21_c54 <= Y_21_c53;
               X_22_c54 <= X_22_c53;
               Y_22_c54 <= Y_22_c53;
            end if;
            if ce_55 = '1' then
               R_1_c55 <= R_1_c54;
               R_2_c55 <= R_2_c54;
               R_3_c55 <= R_3_c54;
               R_4_c55 <= R_4_c54;
               R_5_c55 <= R_5_c54;
               R_6_c55 <= R_6_c54;
               R_7_c55 <= R_7_c54;
               R_8_c55 <= R_8_c54;
               R_9_c55 <= R_9_c54;
               R_10_c55 <= R_10_c54;
               R_11_c55 <= R_11_c54;
               R_12_c55 <= R_12_c54;
               R_13_c55 <= R_13_c54;
               R_14_c55 <= R_14_c54;
               R_15_c55 <= R_15_c54;
               R_16_c55 <= R_16_c54;
               R_17_c55 <= R_17_c54;
               R_18_c55 <= R_18_c54;
               R_19_c55 <= R_19_c54;
               R_20_c55 <= R_20_c54;
               Cin_21_c55 <= Cin_21_c54;
               X_21_c55 <= X_21_c54;
               Y_21_c55 <= Y_21_c54;
               X_22_c55 <= X_22_c54;
               Y_22_c55 <= Y_22_c54;
            end if;
            if ce_56 = '1' then
               R_1_c56 <= R_1_c55;
               R_2_c56 <= R_2_c55;
               R_3_c56 <= R_3_c55;
               R_4_c56 <= R_4_c55;
               R_5_c56 <= R_5_c55;
               R_6_c56 <= R_6_c55;
               R_7_c56 <= R_7_c55;
               R_8_c56 <= R_8_c55;
               R_9_c56 <= R_9_c55;
               R_10_c56 <= R_10_c55;
               R_11_c56 <= R_11_c55;
               R_12_c56 <= R_12_c55;
               R_13_c56 <= R_13_c55;
               R_14_c56 <= R_14_c55;
               R_15_c56 <= R_15_c55;
               R_16_c56 <= R_16_c55;
               R_17_c56 <= R_17_c55;
               R_18_c56 <= R_18_c55;
               R_19_c56 <= R_19_c55;
               R_20_c56 <= R_20_c55;
               Cin_21_c56 <= Cin_21_c55;
               X_21_c56 <= X_21_c55;
               Y_21_c56 <= Y_21_c55;
               X_22_c56 <= X_22_c55;
               Y_22_c56 <= Y_22_c55;
            end if;
         end if;
      end process;
   Cin_1_c34 <= Cin;
   X_1_c33 <= '0' & X(2 downto 0);
   Y_1_c0 <= '0' & Y(2 downto 0);
   S_1_c35 <= X_1_c35 + Y_1_c35 + Cin_1_c35;
   R_1_c35 <= S_1_c35(2 downto 0);
   Cin_2_c35 <= S_1_c35(3);
   X_2_c33 <= '0' & X(5 downto 3);
   Y_2_c0 <= '0' & Y(5 downto 3);
   S_2_c36 <= X_2_c36 + Y_2_c36 + Cin_2_c36;
   R_2_c36 <= S_2_c36(2 downto 0);
   Cin_3_c36 <= S_2_c36(3);
   X_3_c33 <= '0' & X(8 downto 6);
   Y_3_c0 <= '0' & Y(8 downto 6);
   S_3_c37 <= X_3_c37 + Y_3_c37 + Cin_3_c37;
   R_3_c37 <= S_3_c37(2 downto 0);
   Cin_4_c37 <= S_3_c37(3);
   X_4_c33 <= '0' & X(11 downto 9);
   Y_4_c0 <= '0' & Y(11 downto 9);
   S_4_c38 <= X_4_c38 + Y_4_c38 + Cin_4_c38;
   R_4_c38 <= S_4_c38(2 downto 0);
   Cin_5_c38 <= S_4_c38(3);
   X_5_c33 <= '0' & X(14 downto 12);
   Y_5_c0 <= '0' & Y(14 downto 12);
   S_5_c39 <= X_5_c39 + Y_5_c39 + Cin_5_c39;
   R_5_c39 <= S_5_c39(2 downto 0);
   Cin_6_c39 <= S_5_c39(3);
   X_6_c33 <= '0' & X(17 downto 15);
   Y_6_c0 <= '0' & Y(17 downto 15);
   S_6_c40 <= X_6_c40 + Y_6_c40 + Cin_6_c40;
   R_6_c40 <= S_6_c40(2 downto 0);
   Cin_7_c40 <= S_6_c40(3);
   X_7_c33 <= '0' & X(20 downto 18);
   Y_7_c0 <= '0' & Y(20 downto 18);
   S_7_c41 <= X_7_c41 + Y_7_c41 + Cin_7_c41;
   R_7_c41 <= S_7_c41(2 downto 0);
   Cin_8_c41 <= S_7_c41(3);
   X_8_c33 <= '0' & X(23 downto 21);
   Y_8_c0 <= '0' & Y(23 downto 21);
   S_8_c42 <= X_8_c42 + Y_8_c42 + Cin_8_c42;
   R_8_c42 <= S_8_c42(2 downto 0);
   Cin_9_c42 <= S_8_c42(3);
   X_9_c33 <= '0' & X(26 downto 24);
   Y_9_c0 <= '0' & Y(26 downto 24);
   S_9_c43 <= X_9_c43 + Y_9_c43 + Cin_9_c43;
   R_9_c43 <= S_9_c43(2 downto 0);
   Cin_10_c43 <= S_9_c43(3);
   X_10_c33 <= '0' & X(29 downto 27);
   Y_10_c0 <= '0' & Y(29 downto 27);
   S_10_c44 <= X_10_c44 + Y_10_c44 + Cin_10_c44;
   R_10_c44 <= S_10_c44(2 downto 0);
   Cin_11_c44 <= S_10_c44(3);
   X_11_c33 <= '0' & X(32 downto 30);
   Y_11_c0 <= '0' & Y(32 downto 30);
   S_11_c45 <= X_11_c45 + Y_11_c45 + Cin_11_c45;
   R_11_c45 <= S_11_c45(2 downto 0);
   Cin_12_c45 <= S_11_c45(3);
   X_12_c33 <= '0' & X(35 downto 33);
   Y_12_c0 <= '0' & Y(35 downto 33);
   S_12_c46 <= X_12_c46 + Y_12_c46 + Cin_12_c46;
   R_12_c46 <= S_12_c46(2 downto 0);
   Cin_13_c46 <= S_12_c46(3);
   X_13_c33 <= '0' & X(38 downto 36);
   Y_13_c0 <= '0' & Y(38 downto 36);
   S_13_c47 <= X_13_c47 + Y_13_c47 + Cin_13_c47;
   R_13_c47 <= S_13_c47(2 downto 0);
   Cin_14_c47 <= S_13_c47(3);
   X_14_c33 <= '0' & X(41 downto 39);
   Y_14_c0 <= '0' & Y(41 downto 39);
   S_14_c48 <= X_14_c48 + Y_14_c48 + Cin_14_c48;
   R_14_c48 <= S_14_c48(2 downto 0);
   Cin_15_c48 <= S_14_c48(3);
   X_15_c33 <= '0' & X(44 downto 42);
   Y_15_c0 <= '0' & Y(44 downto 42);
   S_15_c49 <= X_15_c49 + Y_15_c49 + Cin_15_c49;
   R_15_c49 <= S_15_c49(2 downto 0);
   Cin_16_c49 <= S_15_c49(3);
   X_16_c33 <= '0' & X(47 downto 45);
   Y_16_c0 <= '0' & Y(47 downto 45);
   S_16_c50 <= X_16_c50 + Y_16_c50 + Cin_16_c50;
   R_16_c50 <= S_16_c50(2 downto 0);
   Cin_17_c50 <= S_16_c50(3);
   X_17_c33 <= '0' & X(50 downto 48);
   Y_17_c0 <= '0' & Y(50 downto 48);
   S_17_c51 <= X_17_c51 + Y_17_c51 + Cin_17_c51;
   R_17_c51 <= S_17_c51(2 downto 0);
   Cin_18_c51 <= S_17_c51(3);
   X_18_c33 <= '0' & X(53 downto 51);
   Y_18_c0 <= '0' & Y(53 downto 51);
   S_18_c52 <= X_18_c52 + Y_18_c52 + Cin_18_c52;
   R_18_c52 <= S_18_c52(2 downto 0);
   Cin_19_c52 <= S_18_c52(3);
   X_19_c33 <= '0' & X(56 downto 54);
   Y_19_c0 <= '0' & Y(56 downto 54);
   S_19_c53 <= X_19_c53 + Y_19_c53 + Cin_19_c53;
   R_19_c53 <= S_19_c53(2 downto 0);
   Cin_20_c53 <= S_19_c53(3);
   X_20_c33 <= '0' & X(59 downto 57);
   Y_20_c0 <= '0' & Y(59 downto 57);
   S_20_c54 <= X_20_c54 + Y_20_c54 + Cin_20_c54;
   R_20_c54 <= S_20_c54(2 downto 0);
   Cin_21_c54 <= S_20_c54(3);
   X_21_c33 <= '0' & X(62 downto 60);
   Y_21_c0 <= '0' & Y(62 downto 60);
   S_21_c56 <= X_21_c56 + Y_21_c56 + Cin_21_c56;
   R_21_c56 <= S_21_c56(2 downto 0);
   Cin_22_c56 <= S_21_c56(3);
   X_22_c33 <= '0' & X(64 downto 63);
   Y_22_c0 <= '0' & Y(64 downto 63);
   S_22_c56 <= X_22_c56 + Y_22_c56 + Cin_22_c56;
   R_22_c56 <= S_22_c56(1 downto 0);
   R <= R_22_c56 & R_21_c56 & R_20_c56 & R_19_c56 & R_18_c56 & R_17_c56 & R_16_c56 & R_15_c56 & R_14_c56 & R_13_c56 & R_12_c56 & R_11_c56 & R_10_c56 & R_9_c56 & R_8_c56 & R_7_c56 & R_6_c56 & R_5_c56 & R_4_c56 & R_3_c56 & R_2_c56 & R_1_c56 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_11_52_uid2_Freq800_uid3)
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier is
   component IntMultiplier_53x53_106_Freq800_uid5 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component IntAdder_65_Freq800_uid975 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3, sign_c4, sign_c5, sign_c6, sign_c7, sign_c8, sign_c9, sign_c10, sign_c11, sign_c12, sign_c13, sign_c14, sign_c15, sign_c16, sign_c17, sign_c18, sign_c19, sign_c20, sign_c21, sign_c22, sign_c23, sign_c24, sign_c25, sign_c26, sign_c27, sign_c28, sign_c29, sign_c30, sign_c31, sign_c32, sign_c33, sign_c34, sign_c35, sign_c36, sign_c37, sign_c38, sign_c39, sign_c40, sign_c41, sign_c42, sign_c43, sign_c44, sign_c45, sign_c46, sign_c47, sign_c48, sign_c49, sign_c50, sign_c51, sign_c52, sign_c53, sign_c54, sign_c55, sign_c56 :  std_logic;
signal expX_c0, expX_c1 :  std_logic_vector(10 downto 0);
signal expY_c0, expY_c1 :  std_logic_vector(10 downto 0);
signal expSumPreSub_c1, expSumPreSub_c2 :  std_logic_vector(12 downto 0);
signal bias_c0, bias_c1, bias_c2 :  std_logic_vector(12 downto 0);
signal expSum_c2, expSum_c3, expSum_c4, expSum_c5, expSum_c6, expSum_c7, expSum_c8, expSum_c9, expSum_c10, expSum_c11, expSum_c12, expSum_c13, expSum_c14, expSum_c15, expSum_c16, expSum_c17, expSum_c18, expSum_c19, expSum_c20, expSum_c21, expSum_c22, expSum_c23, expSum_c24, expSum_c25, expSum_c26, expSum_c27, expSum_c28, expSum_c29, expSum_c30, expSum_c31, expSum_c32, expSum_c33 :  std_logic_vector(12 downto 0);
signal sigX_c0 :  std_logic_vector(52 downto 0);
signal sigY_c0 :  std_logic_vector(52 downto 0);
signal sigProd_c33 :  std_logic_vector(105 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3, exc_c4, exc_c5, exc_c6, exc_c7, exc_c8, exc_c9, exc_c10, exc_c11, exc_c12, exc_c13, exc_c14, exc_c15, exc_c16, exc_c17, exc_c18, exc_c19, exc_c20, exc_c21, exc_c22, exc_c23, exc_c24, exc_c25, exc_c26, exc_c27, exc_c28, exc_c29, exc_c30, exc_c31, exc_c32, exc_c33, exc_c34, exc_c35, exc_c36, exc_c37, exc_c38, exc_c39, exc_c40, exc_c41, exc_c42, exc_c43, exc_c44, exc_c45, exc_c46, exc_c47, exc_c48, exc_c49, exc_c50, exc_c51, exc_c52, exc_c53, exc_c54, exc_c55, exc_c56 :  std_logic_vector(1 downto 0);
signal norm_c33 :  std_logic;
signal expPostNorm_c33 :  std_logic_vector(12 downto 0);
signal sigProdExt_c33, sigProdExt_c34 :  std_logic_vector(105 downto 0);
signal expSig_c33 :  std_logic_vector(64 downto 0);
signal sticky_c33, sticky_c34 :  std_logic;
signal guard_c34 :  std_logic;
signal round_c34 :  std_logic;
signal expSigPostRound_c56 :  std_logic_vector(64 downto 0);
signal excPostNorm_c56 :  std_logic_vector(1 downto 0);
signal finalExc_c56 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expX_c1 <= expX_c0;
               expY_c1 <= expY_c0;
               bias_c1 <= bias_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSumPreSub_c2 <= expSumPreSub_c1;
               bias_c2 <= bias_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               expSum_c3 <= expSum_c2;
               exc_c3 <= exc_c2;
            end if;
            if ce_4 = '1' then
               sign_c4 <= sign_c3;
               expSum_c4 <= expSum_c3;
               exc_c4 <= exc_c3;
            end if;
            if ce_5 = '1' then
               sign_c5 <= sign_c4;
               expSum_c5 <= expSum_c4;
               exc_c5 <= exc_c4;
            end if;
            if ce_6 = '1' then
               sign_c6 <= sign_c5;
               expSum_c6 <= expSum_c5;
               exc_c6 <= exc_c5;
            end if;
            if ce_7 = '1' then
               sign_c7 <= sign_c6;
               expSum_c7 <= expSum_c6;
               exc_c7 <= exc_c6;
            end if;
            if ce_8 = '1' then
               sign_c8 <= sign_c7;
               expSum_c8 <= expSum_c7;
               exc_c8 <= exc_c7;
            end if;
            if ce_9 = '1' then
               sign_c9 <= sign_c8;
               expSum_c9 <= expSum_c8;
               exc_c9 <= exc_c8;
            end if;
            if ce_10 = '1' then
               sign_c10 <= sign_c9;
               expSum_c10 <= expSum_c9;
               exc_c10 <= exc_c9;
            end if;
            if ce_11 = '1' then
               sign_c11 <= sign_c10;
               expSum_c11 <= expSum_c10;
               exc_c11 <= exc_c10;
            end if;
            if ce_12 = '1' then
               sign_c12 <= sign_c11;
               expSum_c12 <= expSum_c11;
               exc_c12 <= exc_c11;
            end if;
            if ce_13 = '1' then
               sign_c13 <= sign_c12;
               expSum_c13 <= expSum_c12;
               exc_c13 <= exc_c12;
            end if;
            if ce_14 = '1' then
               sign_c14 <= sign_c13;
               expSum_c14 <= expSum_c13;
               exc_c14 <= exc_c13;
            end if;
            if ce_15 = '1' then
               sign_c15 <= sign_c14;
               expSum_c15 <= expSum_c14;
               exc_c15 <= exc_c14;
            end if;
            if ce_16 = '1' then
               sign_c16 <= sign_c15;
               expSum_c16 <= expSum_c15;
               exc_c16 <= exc_c15;
            end if;
            if ce_17 = '1' then
               sign_c17 <= sign_c16;
               expSum_c17 <= expSum_c16;
               exc_c17 <= exc_c16;
            end if;
            if ce_18 = '1' then
               sign_c18 <= sign_c17;
               expSum_c18 <= expSum_c17;
               exc_c18 <= exc_c17;
            end if;
            if ce_19 = '1' then
               sign_c19 <= sign_c18;
               expSum_c19 <= expSum_c18;
               exc_c19 <= exc_c18;
            end if;
            if ce_20 = '1' then
               sign_c20 <= sign_c19;
               expSum_c20 <= expSum_c19;
               exc_c20 <= exc_c19;
            end if;
            if ce_21 = '1' then
               sign_c21 <= sign_c20;
               expSum_c21 <= expSum_c20;
               exc_c21 <= exc_c20;
            end if;
            if ce_22 = '1' then
               sign_c22 <= sign_c21;
               expSum_c22 <= expSum_c21;
               exc_c22 <= exc_c21;
            end if;
            if ce_23 = '1' then
               sign_c23 <= sign_c22;
               expSum_c23 <= expSum_c22;
               exc_c23 <= exc_c22;
            end if;
            if ce_24 = '1' then
               sign_c24 <= sign_c23;
               expSum_c24 <= expSum_c23;
               exc_c24 <= exc_c23;
            end if;
            if ce_25 = '1' then
               sign_c25 <= sign_c24;
               expSum_c25 <= expSum_c24;
               exc_c25 <= exc_c24;
            end if;
            if ce_26 = '1' then
               sign_c26 <= sign_c25;
               expSum_c26 <= expSum_c25;
               exc_c26 <= exc_c25;
            end if;
            if ce_27 = '1' then
               sign_c27 <= sign_c26;
               expSum_c27 <= expSum_c26;
               exc_c27 <= exc_c26;
            end if;
            if ce_28 = '1' then
               sign_c28 <= sign_c27;
               expSum_c28 <= expSum_c27;
               exc_c28 <= exc_c27;
            end if;
            if ce_29 = '1' then
               sign_c29 <= sign_c28;
               expSum_c29 <= expSum_c28;
               exc_c29 <= exc_c28;
            end if;
            if ce_30 = '1' then
               sign_c30 <= sign_c29;
               expSum_c30 <= expSum_c29;
               exc_c30 <= exc_c29;
            end if;
            if ce_31 = '1' then
               sign_c31 <= sign_c30;
               expSum_c31 <= expSum_c30;
               exc_c31 <= exc_c30;
            end if;
            if ce_32 = '1' then
               sign_c32 <= sign_c31;
               expSum_c32 <= expSum_c31;
               exc_c32 <= exc_c31;
            end if;
            if ce_33 = '1' then
               sign_c33 <= sign_c32;
               expSum_c33 <= expSum_c32;
               exc_c33 <= exc_c32;
            end if;
            if ce_34 = '1' then
               sign_c34 <= sign_c33;
               exc_c34 <= exc_c33;
               sigProdExt_c34 <= sigProdExt_c33;
               sticky_c34 <= sticky_c33;
            end if;
            if ce_35 = '1' then
               sign_c35 <= sign_c34;
               exc_c35 <= exc_c34;
            end if;
            if ce_36 = '1' then
               sign_c36 <= sign_c35;
               exc_c36 <= exc_c35;
            end if;
            if ce_37 = '1' then
               sign_c37 <= sign_c36;
               exc_c37 <= exc_c36;
            end if;
            if ce_38 = '1' then
               sign_c38 <= sign_c37;
               exc_c38 <= exc_c37;
            end if;
            if ce_39 = '1' then
               sign_c39 <= sign_c38;
               exc_c39 <= exc_c38;
            end if;
            if ce_40 = '1' then
               sign_c40 <= sign_c39;
               exc_c40 <= exc_c39;
            end if;
            if ce_41 = '1' then
               sign_c41 <= sign_c40;
               exc_c41 <= exc_c40;
            end if;
            if ce_42 = '1' then
               sign_c42 <= sign_c41;
               exc_c42 <= exc_c41;
            end if;
            if ce_43 = '1' then
               sign_c43 <= sign_c42;
               exc_c43 <= exc_c42;
            end if;
            if ce_44 = '1' then
               sign_c44 <= sign_c43;
               exc_c44 <= exc_c43;
            end if;
            if ce_45 = '1' then
               sign_c45 <= sign_c44;
               exc_c45 <= exc_c44;
            end if;
            if ce_46 = '1' then
               sign_c46 <= sign_c45;
               exc_c46 <= exc_c45;
            end if;
            if ce_47 = '1' then
               sign_c47 <= sign_c46;
               exc_c47 <= exc_c46;
            end if;
            if ce_48 = '1' then
               sign_c48 <= sign_c47;
               exc_c48 <= exc_c47;
            end if;
            if ce_49 = '1' then
               sign_c49 <= sign_c48;
               exc_c49 <= exc_c48;
            end if;
            if ce_50 = '1' then
               sign_c50 <= sign_c49;
               exc_c50 <= exc_c49;
            end if;
            if ce_51 = '1' then
               sign_c51 <= sign_c50;
               exc_c51 <= exc_c50;
            end if;
            if ce_52 = '1' then
               sign_c52 <= sign_c51;
               exc_c52 <= exc_c51;
            end if;
            if ce_53 = '1' then
               sign_c53 <= sign_c52;
               exc_c53 <= exc_c52;
            end if;
            if ce_54 = '1' then
               sign_c54 <= sign_c53;
               exc_c54 <= exc_c53;
            end if;
            if ce_55 = '1' then
               sign_c55 <= sign_c54;
               exc_c55 <= exc_c54;
            end if;
            if ce_56 = '1' then
               sign_c56 <= sign_c55;
               exc_c56 <= exc_c55;
            end if;
         end if;
      end process;
   sign_c0 <= X(63) xor Y(63);
   expX_c0 <= X(62 downto 52);
   expY_c0 <= Y(62 downto 52);
   expSumPreSub_c1 <= ("00" & expX_c1) + ("00" & expY_c1);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(1023,13);
   expSum_c2 <= expSumPreSub_c2 - bias_c2;
   sigX_c0 <= "1" & X(51 downto 0);
   sigY_c0 <= "1" & Y(51 downto 0);
   SignificandMultiplication: IntMultiplier_53x53_106_Freq800_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c33);
   excSel_c0 <= X(65 downto 64) & Y(65 downto 64);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c33 <= sigProd_c33(105);
   -- exponent update
   expPostNorm_c33 <= expSum_c33 + ("000000000000" & norm_c33);
   -- significand normalization shift
   sigProdExt_c33 <= sigProd_c33(104 downto 0) & "0" when norm_c33='1' else
                         sigProd_c33(103 downto 0) & "00";
   expSig_c33 <= expPostNorm_c33 & sigProdExt_c33(105 downto 54);
   sticky_c33 <= sigProdExt_c33(53);
   guard_c34 <= '0' when sigProdExt_c34(52 downto 0)="00000000000000000000000000000000000000000000000000000" else '1';
   round_c34 <= sticky_c34 and ( (guard_c34 and not(sigProdExt_c34(54))) or (sigProdExt_c34(54) ))  ;
   RoundingAdder: IntAdder_65_Freq800_uid975
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 ce_51=> ce_51,
                 ce_52=> ce_52,
                 ce_53=> ce_53,
                 ce_54=> ce_54,
                 ce_55=> ce_55,
                 ce_56=> ce_56,
                 Cin => round_c34,
                 X => expSig_c33,
                 Y => "00000000000000000000000000000000000000000000000000000000000000000",
                 R => expSigPostRound_c56);
   with expSigPostRound_c56(64 downto 63)  select 
   excPostNorm_c56 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c56  select  
   finalExc_c56 <= exc_c56 when  "11"|"10"|"00",
                       excPostNorm_c56 when others; 
   R <= finalExc_c56 & sign_c56 & expSigPostRound_c56(62 downto 0);
end architecture;



